VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2250.000 BY 840.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END clock
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 836.000 2.210 840.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 836.000 5.890 840.000 ;
    END
  END core_rstn
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END flash_clk
  PIN flash_clk_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 0.000 1081.830 4.000 ;
    END
  END flash_clk_ieb
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END flash_csb
  PIN flash_csb_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END flash_csb_ieb
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.510 0.000 1254.790 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 0.000 1341.270 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.470 0.000 1427.750 4.000 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.850 0.000 1774.130 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.330 0.000 1860.610 4.000 ;
    END
  END flash_io1_oeb
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END flash_io2_oeb
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END gpio_outenb_pad
  PIN jtag_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 319.640 2250.000 320.240 ;
    END
  END jtag_out
  PIN jtag_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 329.160 2250.000 329.760 ;
    END
  END jtag_outenb
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 836.000 13.250 840.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 836.000 1523.430 840.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.870 836.000 1538.150 840.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.050 836.000 1553.330 840.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 836.000 1568.510 840.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.410 836.000 1583.690 840.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.590 836.000 1598.870 840.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 836.000 1614.050 840.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 836.000 1628.770 840.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 836.000 1643.950 840.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 836.000 1659.130 840.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 836.000 164.130 840.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.030 836.000 1674.310 840.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 836.000 1689.490 840.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 836.000 1704.670 840.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.110 836.000 1719.390 840.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.290 836.000 1734.570 840.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.470 836.000 1749.750 840.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 836.000 1764.930 840.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 836.000 1780.110 840.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.010 836.000 1795.290 840.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 836.000 1810.010 840.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 836.000 179.310 840.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.910 836.000 1825.190 840.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.090 836.000 1840.370 840.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.270 836.000 1855.550 840.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.450 836.000 1870.730 840.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.170 836.000 1885.450 840.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.350 836.000 1900.630 840.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.530 836.000 1915.810 840.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.710 836.000 1930.990 840.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 836.000 194.490 840.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 836.000 209.670 840.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 836.000 224.850 840.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 836.000 240.030 840.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 836.000 254.750 840.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 836.000 269.930 840.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 836.000 285.110 840.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 836.000 300.290 840.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 836.000 28.430 840.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 836.000 315.470 840.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 836.000 330.190 840.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 836.000 345.370 840.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 836.000 360.550 840.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 836.000 375.730 840.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 836.000 390.910 840.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 836.000 406.090 840.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 836.000 420.810 840.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 836.000 435.990 840.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 836.000 451.170 840.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 836.000 43.610 840.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 836.000 466.350 840.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 836.000 481.530 840.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 836.000 496.710 840.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 836.000 511.430 840.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 836.000 526.610 840.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 836.000 541.790 840.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 836.000 556.970 840.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 836.000 572.150 840.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 836.000 586.870 840.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 836.000 602.050 840.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 836.000 58.790 840.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 836.000 617.230 840.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 836.000 632.410 840.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 836.000 647.590 840.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 836.000 662.770 840.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 836.000 677.490 840.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 836.000 692.670 840.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 836.000 707.850 840.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 836.000 723.030 840.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 836.000 738.210 840.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 836.000 753.390 840.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 836.000 73.510 840.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 836.000 768.110 840.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 836.000 783.290 840.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 836.000 798.470 840.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 836.000 813.650 840.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 836.000 828.830 840.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 836.000 844.010 840.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 836.000 858.730 840.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 836.000 873.910 840.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 836.000 889.090 840.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 836.000 904.270 840.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 836.000 88.690 840.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 836.000 919.450 840.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 836.000 934.170 840.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 836.000 949.350 840.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 836.000 964.530 840.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 836.000 979.710 840.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 836.000 994.890 840.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 836.000 1010.070 840.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 836.000 1024.790 840.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 836.000 1039.970 840.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 836.000 1055.150 840.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 836.000 103.870 840.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 836.000 1070.330 840.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 836.000 1085.510 840.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.410 836.000 1100.690 840.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 836.000 1115.410 840.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 836.000 1130.590 840.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 836.000 1145.770 840.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 836.000 1160.950 840.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 836.000 1176.130 840.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 836.000 1191.310 840.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 836.000 1206.030 840.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 836.000 119.050 840.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.930 836.000 1221.210 840.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.110 836.000 1236.390 840.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.290 836.000 1251.570 840.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.470 836.000 1266.750 840.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.190 836.000 1281.470 840.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.370 836.000 1296.650 840.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 836.000 1311.830 840.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 836.000 1327.010 840.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 836.000 1342.190 840.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.090 836.000 1357.370 840.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 836.000 134.230 840.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 836.000 1372.090 840.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 836.000 1387.270 840.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.170 836.000 1402.450 840.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 836.000 1417.630 840.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 836.000 1432.810 840.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 836.000 1447.990 840.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 836.000 1462.710 840.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 836.000 1477.890 840.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 836.000 1493.070 840.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.970 836.000 1508.250 840.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 836.000 149.410 840.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 836.000 16.930 840.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 836.000 1527.110 840.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.010 836.000 1542.290 840.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 836.000 1557.470 840.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 836.000 1572.190 840.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 836.000 1587.370 840.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 836.000 1602.550 840.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 836.000 1617.730 840.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 836.000 1632.910 840.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.350 836.000 1647.630 840.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.530 836.000 1662.810 840.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 836.000 168.270 840.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 836.000 1677.990 840.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.890 836.000 1693.170 840.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.070 836.000 1708.350 840.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.250 836.000 1723.530 840.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 836.000 1738.250 840.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1753.150 836.000 1753.430 840.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.330 836.000 1768.610 840.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 836.000 1783.790 840.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.690 836.000 1798.970 840.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.870 836.000 1814.150 840.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 836.000 182.990 840.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.590 836.000 1828.870 840.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.770 836.000 1844.050 840.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.950 836.000 1859.230 840.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 836.000 1874.410 840.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.310 836.000 1889.590 840.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.490 836.000 1904.770 840.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 836.000 1919.490 840.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.390 836.000 1934.670 840.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 836.000 198.170 840.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 836.000 213.350 840.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 836.000 228.530 840.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 836.000 243.710 840.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 836.000 258.890 840.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 836.000 273.610 840.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 836.000 288.790 840.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 836.000 303.970 840.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 836.000 32.110 840.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 836.000 319.150 840.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 836.000 334.330 840.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 836.000 349.050 840.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 836.000 364.230 840.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 836.000 379.410 840.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 836.000 394.590 840.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 836.000 409.770 840.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 836.000 424.950 840.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 836.000 439.670 840.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 836.000 454.850 840.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 836.000 47.290 840.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 836.000 470.030 840.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 836.000 485.210 840.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 836.000 500.390 840.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 836.000 515.570 840.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 836.000 530.290 840.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 836.000 545.470 840.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 836.000 560.650 840.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 836.000 575.830 840.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 836.000 591.010 840.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 836.000 606.190 840.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 836.000 62.470 840.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 836.000 620.910 840.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 836.000 636.090 840.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 836.000 651.270 840.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 836.000 666.450 840.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 836.000 681.630 840.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 836.000 696.350 840.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 836.000 711.530 840.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 836.000 726.710 840.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 836.000 741.890 840.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 836.000 757.070 840.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 836.000 77.650 840.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 836.000 772.250 840.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 836.000 786.970 840.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 836.000 802.150 840.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 836.000 817.330 840.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 836.000 832.510 840.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 836.000 847.690 840.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 836.000 862.870 840.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 836.000 877.590 840.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 836.000 892.770 840.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 836.000 907.950 840.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 836.000 92.370 840.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 836.000 923.130 840.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 836.000 938.310 840.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 836.000 953.490 840.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 836.000 968.210 840.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 836.000 983.390 840.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 836.000 998.570 840.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 836.000 1013.750 840.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 836.000 1028.930 840.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 836.000 1043.650 840.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 836.000 1058.830 840.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 836.000 107.550 840.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 836.000 1074.010 840.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 836.000 1089.190 840.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 836.000 1104.370 840.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 836.000 1119.550 840.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 836.000 1134.270 840.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 836.000 1149.450 840.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 836.000 1164.630 840.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 836.000 1179.810 840.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 836.000 1194.990 840.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.890 836.000 1210.170 840.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 836.000 122.730 840.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.610 836.000 1224.890 840.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 836.000 1240.070 840.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.970 836.000 1255.250 840.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 836.000 1270.430 840.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 836.000 1285.610 840.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 836.000 1300.330 840.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.230 836.000 1315.510 840.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 836.000 1330.690 840.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 836.000 1345.870 840.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 836.000 1361.050 840.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 836.000 137.910 840.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 836.000 1376.230 840.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 836.000 1390.950 840.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 836.000 1406.130 840.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 836.000 1421.310 840.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 836.000 1436.490 840.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 836.000 1451.670 840.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.570 836.000 1466.850 840.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 836.000 1481.570 840.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 836.000 1496.750 840.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 836.000 1511.930 840.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 836.000 153.090 840.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 836.000 21.070 840.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 836.000 1530.790 840.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 836.000 1545.970 840.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 836.000 1561.150 840.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 836.000 1576.330 840.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 836.000 1591.050 840.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 836.000 1606.230 840.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 836.000 1621.410 840.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 836.000 1636.590 840.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 836.000 1651.770 840.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.670 836.000 1666.950 840.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 836.000 171.950 840.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.390 836.000 1681.670 840.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 836.000 1696.850 840.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 836.000 1712.030 840.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.930 836.000 1727.210 840.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 836.000 1742.390 840.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 836.000 1757.110 840.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 836.000 1772.290 840.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 836.000 1787.470 840.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.370 836.000 1802.650 840.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.550 836.000 1817.830 840.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 836.000 187.130 840.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.730 836.000 1833.010 840.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.450 836.000 1847.730 840.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.630 836.000 1862.910 840.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.810 836.000 1878.090 840.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.990 836.000 1893.270 840.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.170 836.000 1908.450 840.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.350 836.000 1923.630 840.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 836.000 1938.350 840.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 836.000 201.850 840.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 836.000 217.030 840.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 836.000 232.210 840.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 836.000 247.390 840.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 836.000 262.570 840.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 836.000 277.750 840.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 836.000 292.470 840.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 836.000 307.650 840.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 836.000 35.790 840.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 836.000 322.830 840.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 836.000 338.010 840.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 836.000 353.190 840.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 836.000 368.370 840.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 836.000 383.090 840.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 836.000 398.270 840.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 836.000 413.450 840.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 836.000 428.630 840.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 836.000 443.810 840.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 836.000 458.530 840.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 836.000 50.970 840.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 836.000 473.710 840.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 836.000 488.890 840.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 836.000 504.070 840.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 836.000 519.250 840.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 836.000 534.430 840.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 836.000 549.150 840.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 836.000 564.330 840.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 836.000 579.510 840.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 836.000 594.690 840.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 836.000 609.870 840.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 836.000 66.150 840.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 836.000 625.050 840.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 836.000 639.770 840.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 836.000 654.950 840.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 836.000 670.130 840.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 836.000 685.310 840.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 836.000 700.490 840.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 836.000 715.670 840.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 836.000 730.390 840.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 836.000 745.570 840.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 836.000 760.750 840.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 836.000 81.330 840.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 836.000 775.930 840.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 836.000 791.110 840.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 836.000 805.830 840.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 836.000 821.010 840.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 836.000 836.190 840.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 836.000 851.370 840.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 836.000 866.550 840.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 836.000 881.730 840.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 836.000 896.450 840.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 836.000 911.630 840.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 836.000 96.510 840.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 836.000 926.810 840.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 836.000 941.990 840.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 836.000 957.170 840.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 836.000 972.350 840.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 836.000 987.070 840.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 836.000 1002.250 840.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 836.000 1017.430 840.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 836.000 1032.610 840.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 836.000 1047.790 840.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 836.000 1062.510 840.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 836.000 111.230 840.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 836.000 1077.690 840.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 836.000 1092.870 840.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 836.000 1108.050 840.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 836.000 1123.230 840.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 836.000 1138.410 840.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 836.000 1153.130 840.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 836.000 1168.310 840.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 836.000 1183.490 840.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 836.000 1198.670 840.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.570 836.000 1213.850 840.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 836.000 126.410 840.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 836.000 1229.030 840.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 836.000 1243.750 840.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 836.000 1258.930 840.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 836.000 1274.110 840.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 836.000 1289.290 840.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 836.000 1304.470 840.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 836.000 1319.650 840.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 836.000 1334.370 840.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 836.000 1349.550 840.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.450 836.000 1364.730 840.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 836.000 141.590 840.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.630 836.000 1379.910 840.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 836.000 1395.090 840.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.530 836.000 1409.810 840.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.710 836.000 1424.990 840.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 836.000 1440.170 840.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 836.000 1455.350 840.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.250 836.000 1470.530 840.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 836.000 1485.710 840.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 836.000 1500.430 840.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 836.000 1515.610 840.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 836.000 156.770 840.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 836.000 24.750 840.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 836.000 1534.470 840.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.370 836.000 1549.650 840.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.550 836.000 1564.830 840.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 836.000 1580.010 840.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 836.000 1595.190 840.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.630 836.000 1609.910 840.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.810 836.000 1625.090 840.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.990 836.000 1640.270 840.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 836.000 1655.450 840.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.350 836.000 1670.630 840.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 836.000 175.630 840.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 836.000 1685.810 840.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 836.000 1700.530 840.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 836.000 1715.710 840.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.610 836.000 1730.890 840.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 836.000 1746.070 840.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 836.000 1761.250 840.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1775.690 836.000 1775.970 840.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.870 836.000 1791.150 840.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.050 836.000 1806.330 840.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.230 836.000 1821.510 840.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 836.000 190.810 840.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.410 836.000 1836.690 840.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 836.000 1851.870 840.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.310 836.000 1866.590 840.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.490 836.000 1881.770 840.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.670 836.000 1896.950 840.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.850 836.000 1912.130 840.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.030 836.000 1927.310 840.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.210 836.000 1942.490 840.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 836.000 205.990 840.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 836.000 220.710 840.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 836.000 235.890 840.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 836.000 251.070 840.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 836.000 266.250 840.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 836.000 281.430 840.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 836.000 296.610 840.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 836.000 311.330 840.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 836.000 39.930 840.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 836.000 326.510 840.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 836.000 341.690 840.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 836.000 356.870 840.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 836.000 372.050 840.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 836.000 387.230 840.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 836.000 401.950 840.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 836.000 417.130 840.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 836.000 432.310 840.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 836.000 447.490 840.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 836.000 462.670 840.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 836.000 54.650 840.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 836.000 477.850 840.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 836.000 492.570 840.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 836.000 507.750 840.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 836.000 522.930 840.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 836.000 538.110 840.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 836.000 553.290 840.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 836.000 568.010 840.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 836.000 583.190 840.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 836.000 598.370 840.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 836.000 613.550 840.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 836.000 69.830 840.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 836.000 628.730 840.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 836.000 643.910 840.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 836.000 658.630 840.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 836.000 673.810 840.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 836.000 688.990 840.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 836.000 704.170 840.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 836.000 719.350 840.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 836.000 734.530 840.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 836.000 749.250 840.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 836.000 764.430 840.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 836.000 85.010 840.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 836.000 779.610 840.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 836.000 794.790 840.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 836.000 809.970 840.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 836.000 824.690 840.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 836.000 839.870 840.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 836.000 855.050 840.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 836.000 870.230 840.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 836.000 885.410 840.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 836.000 900.590 840.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 836.000 915.310 840.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 836.000 100.190 840.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 836.000 930.490 840.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 836.000 945.670 840.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 836.000 960.850 840.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 836.000 976.030 840.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.930 836.000 991.210 840.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 836.000 1005.930 840.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 836.000 1021.110 840.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 836.000 1036.290 840.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 836.000 1051.470 840.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 836.000 1066.650 840.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 836.000 115.370 840.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 836.000 1081.830 840.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 836.000 1096.550 840.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 836.000 1111.730 840.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 836.000 1126.910 840.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 836.000 1142.090 840.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 836.000 1157.270 840.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 836.000 1171.990 840.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 836.000 1187.170 840.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 836.000 1202.350 840.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 836.000 1217.530 840.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 836.000 130.550 840.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 836.000 1232.710 840.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 836.000 1247.890 840.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 836.000 1262.610 840.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 836.000 1277.790 840.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.690 836.000 1292.970 840.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 836.000 1308.150 840.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 836.000 1323.330 840.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 836.000 1338.510 840.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 836.000 1353.230 840.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.130 836.000 1368.410 840.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 836.000 145.270 840.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 836.000 1383.590 840.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.490 836.000 1398.770 840.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 836.000 1413.950 840.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 836.000 1429.130 840.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 836.000 1443.850 840.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 836.000 1459.030 840.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 836.000 1474.210 840.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 836.000 1489.390 840.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 836.000 1504.570 840.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.010 836.000 1519.290 840.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 836.000 160.450 840.000 ;
    END
  END la_output[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 4.800 2250.000 5.400 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 100.000 2250.000 100.600 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 109.520 2250.000 110.120 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 119.040 2250.000 119.640 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 128.560 2250.000 129.160 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 138.080 2250.000 138.680 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 147.600 2250.000 148.200 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 157.120 2250.000 157.720 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 166.640 2250.000 167.240 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 176.160 2250.000 176.760 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 185.680 2250.000 186.280 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 14.320 2250.000 14.920 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 195.200 2250.000 195.800 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 204.720 2250.000 205.320 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 214.240 2250.000 214.840 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 223.760 2250.000 224.360 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 233.280 2250.000 233.880 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 242.800 2250.000 243.400 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 252.320 2250.000 252.920 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 261.840 2250.000 262.440 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 271.360 2250.000 271.960 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 280.880 2250.000 281.480 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 23.840 2250.000 24.440 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 291.080 2250.000 291.680 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 300.600 2250.000 301.200 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 33.360 2250.000 33.960 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 42.880 2250.000 43.480 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 52.400 2250.000 53.000 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 61.920 2250.000 62.520 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 71.440 2250.000 72.040 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 80.960 2250.000 81.560 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 90.480 2250.000 91.080 ;
    END
  END mask_rev[9]
  PIN mgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END mgmt_addr[7]
  PIN mgmt_addr_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END mgmt_addr_ro[0]
  PIN mgmt_addr_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END mgmt_addr_ro[1]
  PIN mgmt_addr_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END mgmt_addr_ro[2]
  PIN mgmt_addr_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END mgmt_addr_ro[3]
  PIN mgmt_addr_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END mgmt_addr_ro[4]
  PIN mgmt_addr_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END mgmt_addr_ro[5]
  PIN mgmt_addr_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END mgmt_addr_ro[6]
  PIN mgmt_addr_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END mgmt_addr_ro[7]
  PIN mgmt_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END mgmt_ena[1]
  PIN mgmt_ena_ro
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END mgmt_ena_ro
  PIN mgmt_in_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 386.280 2250.000 386.880 ;
    END
  END mgmt_in_data[0]
  PIN mgmt_in_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 577.360 2250.000 577.960 ;
    END
  END mgmt_in_data[10]
  PIN mgmt_in_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 596.400 2250.000 597.000 ;
    END
  END mgmt_in_data[11]
  PIN mgmt_in_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 615.440 2250.000 616.040 ;
    END
  END mgmt_in_data[12]
  PIN mgmt_in_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 634.480 2250.000 635.080 ;
    END
  END mgmt_in_data[13]
  PIN mgmt_in_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 653.520 2250.000 654.120 ;
    END
  END mgmt_in_data[14]
  PIN mgmt_in_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 672.560 2250.000 673.160 ;
    END
  END mgmt_in_data[15]
  PIN mgmt_in_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 691.600 2250.000 692.200 ;
    END
  END mgmt_in_data[16]
  PIN mgmt_in_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 710.640 2250.000 711.240 ;
    END
  END mgmt_in_data[17]
  PIN mgmt_in_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 729.680 2250.000 730.280 ;
    END
  END mgmt_in_data[18]
  PIN mgmt_in_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 748.720 2250.000 749.320 ;
    END
  END mgmt_in_data[19]
  PIN mgmt_in_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 405.320 2250.000 405.920 ;
    END
  END mgmt_in_data[1]
  PIN mgmt_in_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 767.760 2250.000 768.360 ;
    END
  END mgmt_in_data[20]
  PIN mgmt_in_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 786.800 2250.000 787.400 ;
    END
  END mgmt_in_data[21]
  PIN mgmt_in_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 805.840 2250.000 806.440 ;
    END
  END mgmt_in_data[22]
  PIN mgmt_in_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 824.880 2250.000 825.480 ;
    END
  END mgmt_in_data[23]
  PIN mgmt_in_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END mgmt_in_data[24]
  PIN mgmt_in_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END mgmt_in_data[25]
  PIN mgmt_in_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mgmt_in_data[26]
  PIN mgmt_in_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END mgmt_in_data[27]
  PIN mgmt_in_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END mgmt_in_data[28]
  PIN mgmt_in_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END mgmt_in_data[29]
  PIN mgmt_in_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 424.360 2250.000 424.960 ;
    END
  END mgmt_in_data[2]
  PIN mgmt_in_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END mgmt_in_data[30]
  PIN mgmt_in_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END mgmt_in_data[31]
  PIN mgmt_in_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END mgmt_in_data[32]
  PIN mgmt_in_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END mgmt_in_data[33]
  PIN mgmt_in_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END mgmt_in_data[34]
  PIN mgmt_in_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END mgmt_in_data[35]
  PIN mgmt_in_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END mgmt_in_data[36]
  PIN mgmt_in_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END mgmt_in_data[37]
  PIN mgmt_in_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 443.400 2250.000 444.000 ;
    END
  END mgmt_in_data[3]
  PIN mgmt_in_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 462.440 2250.000 463.040 ;
    END
  END mgmt_in_data[4]
  PIN mgmt_in_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 481.480 2250.000 482.080 ;
    END
  END mgmt_in_data[5]
  PIN mgmt_in_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 500.520 2250.000 501.120 ;
    END
  END mgmt_in_data[6]
  PIN mgmt_in_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 519.560 2250.000 520.160 ;
    END
  END mgmt_in_data[7]
  PIN mgmt_in_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 538.600 2250.000 539.200 ;
    END
  END mgmt_in_data[8]
  PIN mgmt_in_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 557.640 2250.000 558.240 ;
    END
  END mgmt_in_data[9]
  PIN mgmt_out_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 395.800 2250.000 396.400 ;
    END
  END mgmt_out_data[0]
  PIN mgmt_out_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 586.880 2250.000 587.480 ;
    END
  END mgmt_out_data[10]
  PIN mgmt_out_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 605.920 2250.000 606.520 ;
    END
  END mgmt_out_data[11]
  PIN mgmt_out_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 624.960 2250.000 625.560 ;
    END
  END mgmt_out_data[12]
  PIN mgmt_out_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 644.000 2250.000 644.600 ;
    END
  END mgmt_out_data[13]
  PIN mgmt_out_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 663.040 2250.000 663.640 ;
    END
  END mgmt_out_data[14]
  PIN mgmt_out_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 682.080 2250.000 682.680 ;
    END
  END mgmt_out_data[15]
  PIN mgmt_out_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 701.120 2250.000 701.720 ;
    END
  END mgmt_out_data[16]
  PIN mgmt_out_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 720.160 2250.000 720.760 ;
    END
  END mgmt_out_data[17]
  PIN mgmt_out_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 739.200 2250.000 739.800 ;
    END
  END mgmt_out_data[18]
  PIN mgmt_out_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 758.240 2250.000 758.840 ;
    END
  END mgmt_out_data[19]
  PIN mgmt_out_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 414.840 2250.000 415.440 ;
    END
  END mgmt_out_data[1]
  PIN mgmt_out_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 777.280 2250.000 777.880 ;
    END
  END mgmt_out_data[20]
  PIN mgmt_out_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 796.320 2250.000 796.920 ;
    END
  END mgmt_out_data[21]
  PIN mgmt_out_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 815.360 2250.000 815.960 ;
    END
  END mgmt_out_data[22]
  PIN mgmt_out_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 834.400 2250.000 835.000 ;
    END
  END mgmt_out_data[23]
  PIN mgmt_out_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END mgmt_out_data[24]
  PIN mgmt_out_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.000 4.000 746.600 ;
    END
  END mgmt_out_data[25]
  PIN mgmt_out_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END mgmt_out_data[26]
  PIN mgmt_out_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.960 4.000 761.560 ;
    END
  END mgmt_out_data[27]
  PIN mgmt_out_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END mgmt_out_data[28]
  PIN mgmt_out_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END mgmt_out_data[29]
  PIN mgmt_out_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 433.880 2250.000 434.480 ;
    END
  END mgmt_out_data[2]
  PIN mgmt_out_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.080 4.000 784.680 ;
    END
  END mgmt_out_data[30]
  PIN mgmt_out_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END mgmt_out_data[31]
  PIN mgmt_out_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END mgmt_out_data[32]
  PIN mgmt_out_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END mgmt_out_data[33]
  PIN mgmt_out_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.000 4.000 814.600 ;
    END
  END mgmt_out_data[34]
  PIN mgmt_out_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END mgmt_out_data[35]
  PIN mgmt_out_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END mgmt_out_data[36]
  PIN mgmt_out_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END mgmt_out_data[37]
  PIN mgmt_out_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 452.920 2250.000 453.520 ;
    END
  END mgmt_out_data[3]
  PIN mgmt_out_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 471.960 2250.000 472.560 ;
    END
  END mgmt_out_data[4]
  PIN mgmt_out_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 491.000 2250.000 491.600 ;
    END
  END mgmt_out_data[5]
  PIN mgmt_out_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 510.040 2250.000 510.640 ;
    END
  END mgmt_out_data[6]
  PIN mgmt_out_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 529.080 2250.000 529.680 ;
    END
  END mgmt_out_data[7]
  PIN mgmt_out_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 548.120 2250.000 548.720 ;
    END
  END mgmt_out_data[8]
  PIN mgmt_out_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 567.840 2250.000 568.440 ;
    END
  END mgmt_out_data[9]
  PIN mgmt_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 521.600 4.000 522.200 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_rdata_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END mgmt_rdata_ro[0]
  PIN mgmt_rdata_ro[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END mgmt_rdata_ro[10]
  PIN mgmt_rdata_ro[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END mgmt_rdata_ro[11]
  PIN mgmt_rdata_ro[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END mgmt_rdata_ro[12]
  PIN mgmt_rdata_ro[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END mgmt_rdata_ro[13]
  PIN mgmt_rdata_ro[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END mgmt_rdata_ro[14]
  PIN mgmt_rdata_ro[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END mgmt_rdata_ro[15]
  PIN mgmt_rdata_ro[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END mgmt_rdata_ro[16]
  PIN mgmt_rdata_ro[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END mgmt_rdata_ro[17]
  PIN mgmt_rdata_ro[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mgmt_rdata_ro[18]
  PIN mgmt_rdata_ro[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END mgmt_rdata_ro[19]
  PIN mgmt_rdata_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END mgmt_rdata_ro[1]
  PIN mgmt_rdata_ro[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END mgmt_rdata_ro[20]
  PIN mgmt_rdata_ro[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END mgmt_rdata_ro[21]
  PIN mgmt_rdata_ro[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END mgmt_rdata_ro[22]
  PIN mgmt_rdata_ro[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END mgmt_rdata_ro[23]
  PIN mgmt_rdata_ro[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END mgmt_rdata_ro[24]
  PIN mgmt_rdata_ro[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END mgmt_rdata_ro[25]
  PIN mgmt_rdata_ro[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END mgmt_rdata_ro[26]
  PIN mgmt_rdata_ro[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END mgmt_rdata_ro[27]
  PIN mgmt_rdata_ro[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END mgmt_rdata_ro[28]
  PIN mgmt_rdata_ro[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mgmt_rdata_ro[29]
  PIN mgmt_rdata_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END mgmt_rdata_ro[2]
  PIN mgmt_rdata_ro[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END mgmt_rdata_ro[30]
  PIN mgmt_rdata_ro[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END mgmt_rdata_ro[31]
  PIN mgmt_rdata_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END mgmt_rdata_ro[3]
  PIN mgmt_rdata_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END mgmt_rdata_ro[4]
  PIN mgmt_rdata_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END mgmt_rdata_ro[5]
  PIN mgmt_rdata_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END mgmt_rdata_ro[6]
  PIN mgmt_rdata_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END mgmt_rdata_ro[7]
  PIN mgmt_rdata_ro[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END mgmt_rdata_ro[8]
  PIN mgmt_rdata_ro[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END mgmt_rdata_ro[9]
  PIN mgmt_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END mgmt_wen_mask[7]
  PIN mprj2_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2217.750 836.000 2218.030 840.000 ;
    END
  END mprj2_vcc_pwrgood
  PIN mprj2_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 836.000 2225.390 840.000 ;
    END
  END mprj2_vdd_pwrgood
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.930 836.000 1957.210 840.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.550 836.000 2047.830 840.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.370 836.000 2055.650 840.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.730 836.000 2063.010 840.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 836.000 2070.830 840.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.910 836.000 2078.190 840.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.270 836.000 2085.550 840.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.090 836.000 2093.370 840.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.450 836.000 2100.730 840.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.270 836.000 2108.550 840.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 836.000 2115.910 840.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.430 836.000 1968.710 840.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.990 836.000 2123.270 840.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.810 836.000 2131.090 840.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 836.000 2138.450 840.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.990 836.000 2146.270 840.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.350 836.000 2153.630 840.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.170 836.000 2161.450 840.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.530 836.000 2168.810 840.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.890 836.000 2176.170 840.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.710 836.000 2183.990 840.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.070 836.000 2191.350 840.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.930 836.000 1980.210 840.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.890 836.000 2199.170 840.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.250 836.000 2206.530 840.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.970 836.000 1991.250 840.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.470 836.000 2002.750 840.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.830 836.000 2010.110 840.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.650 836.000 2017.930 840.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.010 836.000 2025.290 840.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2032.830 836.000 2033.110 840.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.190 836.000 2040.470 840.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.890 836.000 1946.170 840.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 836.000 1961.350 840.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.690 836.000 2051.970 840.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.050 836.000 2059.330 840.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.410 836.000 2066.690 840.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2074.230 836.000 2074.510 840.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.590 836.000 2081.870 840.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.410 836.000 2089.690 840.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.770 836.000 2097.050 840.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.130 836.000 2104.410 840.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.950 836.000 2112.230 840.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.310 836.000 2119.590 840.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 836.000 1972.390 840.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.130 836.000 2127.410 840.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.490 836.000 2134.770 840.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.310 836.000 2142.590 840.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.670 836.000 2149.950 840.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.030 836.000 2157.310 840.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.850 836.000 2165.130 840.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.210 836.000 2172.490 840.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 836.000 2180.310 840.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2187.390 836.000 2187.670 840.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.750 836.000 2195.030 840.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 836.000 1983.890 840.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.570 836.000 2202.850 840.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.930 836.000 2210.210 840.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.650 836.000 1994.930 840.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.150 836.000 2006.430 840.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.510 836.000 2013.790 840.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.330 836.000 2021.610 840.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 836.000 2028.970 840.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.510 836.000 2036.790 840.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.870 836.000 2044.150 840.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_io_loader_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 348.200 2250.000 348.800 ;
    END
  END mprj_io_loader_clock
  PIN mprj_io_loader_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 376.760 2250.000 377.360 ;
    END
  END mprj_io_loader_data_1
  PIN mprj_io_loader_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END mprj_io_loader_data_2
  PIN mprj_io_loader_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 338.680 2250.000 339.280 ;
    END
  END mprj_io_loader_resetn
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.750 836.000 1965.030 840.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 836.000 1976.070 840.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.290 836.000 1987.570 840.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.790 836.000 1999.070 840.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.570 836.000 1949.850 840.000 ;
    END
  END mprj_stb_o
  PIN mprj_vcc_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.610 836.000 2213.890 840.000 ;
    END
  END mprj_vcc_pwrgood
  PIN mprj_vdd_pwrgood
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.430 836.000 2221.710 840.000 ;
    END
  END mprj_vdd_pwrgood
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.250 836.000 1953.530 840.000 ;
    END
  END mprj_we_o
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 310.120 2250.000 310.720 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.810 0.000 1947.090 4.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.290 0.000 2033.570 4.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.770 0.000 2120.050 4.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.250 0.000 2206.530 4.000 ;
    END
  END pwr_ctrl_out[3]
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END resetb
  PIN sdo_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 357.720 2250.000 358.320 ;
    END
  END sdo_out
  PIN sdo_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 367.240 2250.000 367.840 ;
    END
  END sdo_outenb
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 836.000 9.570 840.000 ;
    END
  END user_clk
  PIN user_irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 836.000 2229.070 840.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.470 836.000 2232.750 840.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.610 836.000 2236.890 840.000 ;
    END
  END user_irq[2]
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.290 836.000 2240.570 840.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.970 836.000 2244.250 840.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 836.000 2247.930 840.000 ;
    END
  END user_irq_ena[2]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2221.040 10.640 2222.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.040 10.640 2172.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2121.040 10.640 2122.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2071.040 10.640 2072.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2021.040 10.640 2022.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1971.040 821.480 1972.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1921.040 10.640 1922.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1871.040 10.640 1872.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1821.040 10.640 1822.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1771.040 10.640 1772.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1721.040 10.640 1722.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1671.040 10.640 1672.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1621.040 10.640 1622.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 640.760 872.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 640.760 822.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 640.760 772.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 640.760 722.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 640.760 672.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 640.760 622.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 640.760 572.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 640.760 522.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 640.760 472.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 640.760 422.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 640.760 372.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 640.760 322.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 640.760 272.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 640.760 222.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 640.760 172.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 640.760 122.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 827.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1971.040 10.640 1972.640 726.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 106.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 806.490 2244.340 808.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 676.490 2244.340 678.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 546.490 2244.340 548.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 416.490 2244.340 418.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 286.490 2244.340 288.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 156.490 2244.340 158.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2244.340 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2196.040 10.640 2197.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2146.040 10.640 2147.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2096.040 10.640 2097.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2046.040 10.640 2047.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1996.040 821.480 1997.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1946.040 821.480 1947.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1896.040 10.640 1897.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1846.040 10.640 1847.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1796.040 10.640 1797.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1746.040 10.640 1747.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1696.040 10.640 1697.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1646.040 10.640 1647.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1596.040 10.640 1597.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1546.040 10.640 1547.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1496.040 10.640 1497.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1446.040 10.640 1447.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1396.040 10.640 1397.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1346.040 10.640 1347.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1296.040 10.640 1297.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1246.040 10.640 1247.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1196.040 10.640 1197.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 640.760 847.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 640.760 797.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 640.760 747.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 640.760 697.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 640.760 647.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 640.760 597.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 640.760 547.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 640.760 497.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 640.760 447.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 640.760 397.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 640.760 347.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 640.760 297.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 640.760 247.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 640.760 197.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 640.760 147.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 827.120 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1996.040 10.640 1997.640 726.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1946.040 10.640 1947.640 726.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 106.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 741.490 2244.340 743.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 611.490 2244.340 613.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 481.490 2244.340 483.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 351.490 2244.340 353.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 221.490 2244.340 223.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 91.490 2244.340 93.090 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2244.340 836.995 ;
      LAYER met1 ;
        RECT 393.830 840.040 394.150 840.100 ;
        RECT 880.510 840.040 880.830 840.100 ;
        RECT 393.830 840.000 880.830 840.040 ;
        RECT 999.190 840.040 999.510 840.100 ;
        RECT 1384.210 840.040 1384.530 840.100 ;
        RECT 999.190 840.000 1384.530 840.040 ;
        RECT 0.070 5.140 2247.490 840.000 ;
      LAYER met2 ;
        RECT 393.860 840.000 394.120 840.130 ;
        RECT 880.540 840.000 880.800 840.130 ;
        RECT 999.220 840.000 999.480 840.130 ;
        RECT 1384.240 840.000 1384.500 840.130 ;
        RECT 0.090 835.720 1.650 840.000 ;
        RECT 2.490 835.720 5.330 840.000 ;
        RECT 6.170 835.720 9.010 840.000 ;
        RECT 9.850 835.720 12.690 840.000 ;
        RECT 13.530 835.720 16.370 840.000 ;
        RECT 17.210 835.720 20.510 840.000 ;
        RECT 21.350 835.720 24.190 840.000 ;
        RECT 25.030 835.720 27.870 840.000 ;
        RECT 28.710 835.720 31.550 840.000 ;
        RECT 32.390 835.720 35.230 840.000 ;
        RECT 36.070 835.720 39.370 840.000 ;
        RECT 40.210 835.720 43.050 840.000 ;
        RECT 43.890 835.720 46.730 840.000 ;
        RECT 47.570 835.720 50.410 840.000 ;
        RECT 51.250 835.720 54.090 840.000 ;
        RECT 54.930 835.720 58.230 840.000 ;
        RECT 59.070 835.720 61.910 840.000 ;
        RECT 62.750 835.720 65.590 840.000 ;
        RECT 66.430 835.720 69.270 840.000 ;
        RECT 70.110 835.720 72.950 840.000 ;
        RECT 73.790 835.720 77.090 840.000 ;
        RECT 77.930 835.720 80.770 840.000 ;
        RECT 81.610 835.720 84.450 840.000 ;
        RECT 85.290 835.720 88.130 840.000 ;
        RECT 88.970 835.720 91.810 840.000 ;
        RECT 92.650 835.720 95.950 840.000 ;
        RECT 96.790 835.720 99.630 840.000 ;
        RECT 100.470 835.720 103.310 840.000 ;
        RECT 104.150 835.720 106.990 840.000 ;
        RECT 107.830 835.720 110.670 840.000 ;
        RECT 111.510 835.720 114.810 840.000 ;
        RECT 115.650 835.720 118.490 840.000 ;
        RECT 119.330 835.720 122.170 840.000 ;
        RECT 123.010 835.720 125.850 840.000 ;
        RECT 126.690 835.720 129.990 840.000 ;
        RECT 130.830 835.720 133.670 840.000 ;
        RECT 134.510 835.720 137.350 840.000 ;
        RECT 138.190 835.720 141.030 840.000 ;
        RECT 141.870 835.720 144.710 840.000 ;
        RECT 145.550 835.720 148.850 840.000 ;
        RECT 149.690 835.720 152.530 840.000 ;
        RECT 153.370 835.720 156.210 840.000 ;
        RECT 157.050 835.720 159.890 840.000 ;
        RECT 160.730 835.720 163.570 840.000 ;
        RECT 164.410 835.720 167.710 840.000 ;
        RECT 168.550 835.720 171.390 840.000 ;
        RECT 172.230 835.720 175.070 840.000 ;
        RECT 175.910 835.720 178.750 840.000 ;
        RECT 179.590 835.720 182.430 840.000 ;
        RECT 183.270 835.720 186.570 840.000 ;
        RECT 187.410 835.720 190.250 840.000 ;
        RECT 191.090 835.720 193.930 840.000 ;
        RECT 194.770 835.720 197.610 840.000 ;
        RECT 198.450 835.720 201.290 840.000 ;
        RECT 202.130 835.720 205.430 840.000 ;
        RECT 206.270 835.720 209.110 840.000 ;
        RECT 209.950 835.720 212.790 840.000 ;
        RECT 213.630 835.720 216.470 840.000 ;
        RECT 217.310 835.720 220.150 840.000 ;
        RECT 220.990 835.720 224.290 840.000 ;
        RECT 225.130 835.720 227.970 840.000 ;
        RECT 228.810 835.720 231.650 840.000 ;
        RECT 232.490 835.720 235.330 840.000 ;
        RECT 236.170 835.720 239.470 840.000 ;
        RECT 240.310 835.720 243.150 840.000 ;
        RECT 243.990 835.720 246.830 840.000 ;
        RECT 247.670 835.720 250.510 840.000 ;
        RECT 251.350 835.720 254.190 840.000 ;
        RECT 255.030 835.720 258.330 840.000 ;
        RECT 259.170 835.720 262.010 840.000 ;
        RECT 262.850 835.720 265.690 840.000 ;
        RECT 266.530 835.720 269.370 840.000 ;
        RECT 270.210 835.720 273.050 840.000 ;
        RECT 273.890 835.720 277.190 840.000 ;
        RECT 278.030 835.720 280.870 840.000 ;
        RECT 281.710 835.720 284.550 840.000 ;
        RECT 285.390 835.720 288.230 840.000 ;
        RECT 289.070 835.720 291.910 840.000 ;
        RECT 292.750 835.720 296.050 840.000 ;
        RECT 296.890 835.720 299.730 840.000 ;
        RECT 300.570 835.720 303.410 840.000 ;
        RECT 304.250 835.720 307.090 840.000 ;
        RECT 307.930 835.720 310.770 840.000 ;
        RECT 311.610 835.720 314.910 840.000 ;
        RECT 315.750 835.720 318.590 840.000 ;
        RECT 319.430 835.720 322.270 840.000 ;
        RECT 323.110 835.720 325.950 840.000 ;
        RECT 326.790 835.720 329.630 840.000 ;
        RECT 330.470 835.720 333.770 840.000 ;
        RECT 334.610 835.720 337.450 840.000 ;
        RECT 338.290 835.720 341.130 840.000 ;
        RECT 341.970 835.720 344.810 840.000 ;
        RECT 345.650 835.720 348.490 840.000 ;
        RECT 349.330 835.720 352.630 840.000 ;
        RECT 353.470 835.720 356.310 840.000 ;
        RECT 357.150 835.720 359.990 840.000 ;
        RECT 360.830 835.720 363.670 840.000 ;
        RECT 364.510 835.720 367.810 840.000 ;
        RECT 368.650 835.720 371.490 840.000 ;
        RECT 372.330 835.720 375.170 840.000 ;
        RECT 376.010 835.720 378.850 840.000 ;
        RECT 379.690 835.720 382.530 840.000 ;
        RECT 383.370 835.720 386.670 840.000 ;
        RECT 387.510 835.720 390.350 840.000 ;
        RECT 391.190 839.840 394.120 840.000 ;
        RECT 391.190 835.720 394.030 839.840 ;
        RECT 394.870 835.720 397.710 840.000 ;
        RECT 398.550 835.720 401.390 840.000 ;
        RECT 402.230 835.720 405.530 840.000 ;
        RECT 406.370 835.720 409.210 840.000 ;
        RECT 410.050 835.720 412.890 840.000 ;
        RECT 413.730 835.720 416.570 840.000 ;
        RECT 417.410 835.720 420.250 840.000 ;
        RECT 421.090 835.720 424.390 840.000 ;
        RECT 425.230 835.720 428.070 840.000 ;
        RECT 428.910 835.720 431.750 840.000 ;
        RECT 432.590 835.720 435.430 840.000 ;
        RECT 436.270 835.720 439.110 840.000 ;
        RECT 439.950 835.720 443.250 840.000 ;
        RECT 444.090 835.720 446.930 840.000 ;
        RECT 447.770 835.720 450.610 840.000 ;
        RECT 451.450 835.720 454.290 840.000 ;
        RECT 455.130 835.720 457.970 840.000 ;
        RECT 458.810 835.720 462.110 840.000 ;
        RECT 462.950 835.720 465.790 840.000 ;
        RECT 466.630 835.720 469.470 840.000 ;
        RECT 470.310 835.720 473.150 840.000 ;
        RECT 473.990 835.720 477.290 840.000 ;
        RECT 478.130 835.720 480.970 840.000 ;
        RECT 481.810 835.720 484.650 840.000 ;
        RECT 485.490 835.720 488.330 840.000 ;
        RECT 489.170 835.720 492.010 840.000 ;
        RECT 492.850 835.720 496.150 840.000 ;
        RECT 496.990 835.720 499.830 840.000 ;
        RECT 500.670 835.720 503.510 840.000 ;
        RECT 504.350 835.720 507.190 840.000 ;
        RECT 508.030 835.720 510.870 840.000 ;
        RECT 511.710 835.720 515.010 840.000 ;
        RECT 515.850 835.720 518.690 840.000 ;
        RECT 519.530 835.720 522.370 840.000 ;
        RECT 523.210 835.720 526.050 840.000 ;
        RECT 526.890 835.720 529.730 840.000 ;
        RECT 530.570 835.720 533.870 840.000 ;
        RECT 534.710 835.720 537.550 840.000 ;
        RECT 538.390 835.720 541.230 840.000 ;
        RECT 542.070 835.720 544.910 840.000 ;
        RECT 545.750 835.720 548.590 840.000 ;
        RECT 549.430 835.720 552.730 840.000 ;
        RECT 553.570 835.720 556.410 840.000 ;
        RECT 557.250 835.720 560.090 840.000 ;
        RECT 560.930 835.720 563.770 840.000 ;
        RECT 564.610 835.720 567.450 840.000 ;
        RECT 568.290 835.720 571.590 840.000 ;
        RECT 572.430 835.720 575.270 840.000 ;
        RECT 576.110 835.720 578.950 840.000 ;
        RECT 579.790 835.720 582.630 840.000 ;
        RECT 583.470 835.720 586.310 840.000 ;
        RECT 587.150 835.720 590.450 840.000 ;
        RECT 591.290 835.720 594.130 840.000 ;
        RECT 594.970 835.720 597.810 840.000 ;
        RECT 598.650 835.720 601.490 840.000 ;
        RECT 602.330 835.720 605.630 840.000 ;
        RECT 606.470 835.720 609.310 840.000 ;
        RECT 610.150 835.720 612.990 840.000 ;
        RECT 613.830 835.720 616.670 840.000 ;
        RECT 617.510 835.720 620.350 840.000 ;
        RECT 621.190 835.720 624.490 840.000 ;
        RECT 625.330 835.720 628.170 840.000 ;
        RECT 629.010 835.720 631.850 840.000 ;
        RECT 632.690 835.720 635.530 840.000 ;
        RECT 636.370 835.720 639.210 840.000 ;
        RECT 640.050 835.720 643.350 840.000 ;
        RECT 644.190 835.720 647.030 840.000 ;
        RECT 647.870 835.720 650.710 840.000 ;
        RECT 651.550 835.720 654.390 840.000 ;
        RECT 655.230 835.720 658.070 840.000 ;
        RECT 658.910 835.720 662.210 840.000 ;
        RECT 663.050 835.720 665.890 840.000 ;
        RECT 666.730 835.720 669.570 840.000 ;
        RECT 670.410 835.720 673.250 840.000 ;
        RECT 674.090 835.720 676.930 840.000 ;
        RECT 677.770 835.720 681.070 840.000 ;
        RECT 681.910 835.720 684.750 840.000 ;
        RECT 685.590 835.720 688.430 840.000 ;
        RECT 689.270 835.720 692.110 840.000 ;
        RECT 692.950 835.720 695.790 840.000 ;
        RECT 696.630 835.720 699.930 840.000 ;
        RECT 700.770 835.720 703.610 840.000 ;
        RECT 704.450 835.720 707.290 840.000 ;
        RECT 708.130 835.720 710.970 840.000 ;
        RECT 711.810 835.720 715.110 840.000 ;
        RECT 715.950 835.720 718.790 840.000 ;
        RECT 719.630 835.720 722.470 840.000 ;
        RECT 723.310 835.720 726.150 840.000 ;
        RECT 726.990 835.720 729.830 840.000 ;
        RECT 730.670 835.720 733.970 840.000 ;
        RECT 734.810 835.720 737.650 840.000 ;
        RECT 738.490 835.720 741.330 840.000 ;
        RECT 742.170 835.720 745.010 840.000 ;
        RECT 745.850 835.720 748.690 840.000 ;
        RECT 749.530 835.720 752.830 840.000 ;
        RECT 753.670 835.720 756.510 840.000 ;
        RECT 757.350 835.720 760.190 840.000 ;
        RECT 761.030 835.720 763.870 840.000 ;
        RECT 764.710 835.720 767.550 840.000 ;
        RECT 768.390 835.720 771.690 840.000 ;
        RECT 772.530 835.720 775.370 840.000 ;
        RECT 776.210 835.720 779.050 840.000 ;
        RECT 779.890 835.720 782.730 840.000 ;
        RECT 783.570 835.720 786.410 840.000 ;
        RECT 787.250 835.720 790.550 840.000 ;
        RECT 791.390 835.720 794.230 840.000 ;
        RECT 795.070 835.720 797.910 840.000 ;
        RECT 798.750 835.720 801.590 840.000 ;
        RECT 802.430 835.720 805.270 840.000 ;
        RECT 806.110 835.720 809.410 840.000 ;
        RECT 810.250 835.720 813.090 840.000 ;
        RECT 813.930 835.720 816.770 840.000 ;
        RECT 817.610 835.720 820.450 840.000 ;
        RECT 821.290 835.720 824.130 840.000 ;
        RECT 824.970 835.720 828.270 840.000 ;
        RECT 829.110 835.720 831.950 840.000 ;
        RECT 832.790 835.720 835.630 840.000 ;
        RECT 836.470 835.720 839.310 840.000 ;
        RECT 840.150 835.720 843.450 840.000 ;
        RECT 844.290 835.720 847.130 840.000 ;
        RECT 847.970 835.720 850.810 840.000 ;
        RECT 851.650 835.720 854.490 840.000 ;
        RECT 855.330 835.720 858.170 840.000 ;
        RECT 859.010 835.720 862.310 840.000 ;
        RECT 863.150 835.720 865.990 840.000 ;
        RECT 866.830 835.720 869.670 840.000 ;
        RECT 870.510 835.720 873.350 840.000 ;
        RECT 874.190 835.720 877.030 840.000 ;
        RECT 877.870 835.720 881.170 840.000 ;
        RECT 882.010 835.720 884.850 840.000 ;
        RECT 885.690 835.720 888.530 840.000 ;
        RECT 889.370 835.720 892.210 840.000 ;
        RECT 893.050 835.720 895.890 840.000 ;
        RECT 896.730 835.720 900.030 840.000 ;
        RECT 900.870 835.720 903.710 840.000 ;
        RECT 904.550 835.720 907.390 840.000 ;
        RECT 908.230 835.720 911.070 840.000 ;
        RECT 911.910 835.720 914.750 840.000 ;
        RECT 915.590 835.720 918.890 840.000 ;
        RECT 919.730 835.720 922.570 840.000 ;
        RECT 923.410 835.720 926.250 840.000 ;
        RECT 927.090 835.720 929.930 840.000 ;
        RECT 930.770 835.720 933.610 840.000 ;
        RECT 934.450 835.720 937.750 840.000 ;
        RECT 938.590 835.720 941.430 840.000 ;
        RECT 942.270 835.720 945.110 840.000 ;
        RECT 945.950 835.720 948.790 840.000 ;
        RECT 949.630 835.720 952.930 840.000 ;
        RECT 953.770 835.720 956.610 840.000 ;
        RECT 957.450 835.720 960.290 840.000 ;
        RECT 961.130 835.720 963.970 840.000 ;
        RECT 964.810 835.720 967.650 840.000 ;
        RECT 968.490 835.720 971.790 840.000 ;
        RECT 972.630 835.720 975.470 840.000 ;
        RECT 976.310 835.720 979.150 840.000 ;
        RECT 979.990 835.720 982.830 840.000 ;
        RECT 983.670 835.720 986.510 840.000 ;
        RECT 987.350 835.720 990.650 840.000 ;
        RECT 991.490 835.720 994.330 840.000 ;
        RECT 995.170 835.720 998.010 840.000 ;
        RECT 998.850 835.720 1001.690 840.000 ;
        RECT 1002.530 835.720 1005.370 840.000 ;
        RECT 1006.210 835.720 1009.510 840.000 ;
        RECT 1010.350 835.720 1013.190 840.000 ;
        RECT 1014.030 835.720 1016.870 840.000 ;
        RECT 1017.710 835.720 1020.550 840.000 ;
        RECT 1021.390 835.720 1024.230 840.000 ;
        RECT 1025.070 835.720 1028.370 840.000 ;
        RECT 1029.210 835.720 1032.050 840.000 ;
        RECT 1032.890 835.720 1035.730 840.000 ;
        RECT 1036.570 835.720 1039.410 840.000 ;
        RECT 1040.250 835.720 1043.090 840.000 ;
        RECT 1043.930 835.720 1047.230 840.000 ;
        RECT 1048.070 835.720 1050.910 840.000 ;
        RECT 1051.750 835.720 1054.590 840.000 ;
        RECT 1055.430 835.720 1058.270 840.000 ;
        RECT 1059.110 835.720 1061.950 840.000 ;
        RECT 1062.790 835.720 1066.090 840.000 ;
        RECT 1066.930 835.720 1069.770 840.000 ;
        RECT 1070.610 835.720 1073.450 840.000 ;
        RECT 1074.290 835.720 1077.130 840.000 ;
        RECT 1077.970 835.720 1081.270 840.000 ;
        RECT 1082.110 835.720 1084.950 840.000 ;
        RECT 1085.790 835.720 1088.630 840.000 ;
        RECT 1089.470 835.720 1092.310 840.000 ;
        RECT 1093.150 835.720 1095.990 840.000 ;
        RECT 1096.830 835.720 1100.130 840.000 ;
        RECT 1100.970 835.720 1103.810 840.000 ;
        RECT 1104.650 835.720 1107.490 840.000 ;
        RECT 1108.330 835.720 1111.170 840.000 ;
        RECT 1112.010 835.720 1114.850 840.000 ;
        RECT 1115.690 835.720 1118.990 840.000 ;
        RECT 1119.830 835.720 1122.670 840.000 ;
        RECT 1123.510 835.720 1126.350 840.000 ;
        RECT 1127.190 835.720 1130.030 840.000 ;
        RECT 1130.870 835.720 1133.710 840.000 ;
        RECT 1134.550 835.720 1137.850 840.000 ;
        RECT 1138.690 835.720 1141.530 840.000 ;
        RECT 1142.370 835.720 1145.210 840.000 ;
        RECT 1146.050 835.720 1148.890 840.000 ;
        RECT 1149.730 835.720 1152.570 840.000 ;
        RECT 1153.410 835.720 1156.710 840.000 ;
        RECT 1157.550 835.720 1160.390 840.000 ;
        RECT 1161.230 835.720 1164.070 840.000 ;
        RECT 1164.910 835.720 1167.750 840.000 ;
        RECT 1168.590 835.720 1171.430 840.000 ;
        RECT 1172.270 835.720 1175.570 840.000 ;
        RECT 1176.410 835.720 1179.250 840.000 ;
        RECT 1180.090 835.720 1182.930 840.000 ;
        RECT 1183.770 835.720 1186.610 840.000 ;
        RECT 1187.450 835.720 1190.750 840.000 ;
        RECT 1191.590 835.720 1194.430 840.000 ;
        RECT 1195.270 835.720 1198.110 840.000 ;
        RECT 1198.950 835.720 1201.790 840.000 ;
        RECT 1202.630 835.720 1205.470 840.000 ;
        RECT 1206.310 835.720 1209.610 840.000 ;
        RECT 1210.450 835.720 1213.290 840.000 ;
        RECT 1214.130 835.720 1216.970 840.000 ;
        RECT 1217.810 835.720 1220.650 840.000 ;
        RECT 1221.490 835.720 1224.330 840.000 ;
        RECT 1225.170 835.720 1228.470 840.000 ;
        RECT 1229.310 835.720 1232.150 840.000 ;
        RECT 1232.990 835.720 1235.830 840.000 ;
        RECT 1236.670 835.720 1239.510 840.000 ;
        RECT 1240.350 835.720 1243.190 840.000 ;
        RECT 1244.030 835.720 1247.330 840.000 ;
        RECT 1248.170 835.720 1251.010 840.000 ;
        RECT 1251.850 835.720 1254.690 840.000 ;
        RECT 1255.530 835.720 1258.370 840.000 ;
        RECT 1259.210 835.720 1262.050 840.000 ;
        RECT 1262.890 835.720 1266.190 840.000 ;
        RECT 1267.030 835.720 1269.870 840.000 ;
        RECT 1270.710 835.720 1273.550 840.000 ;
        RECT 1274.390 835.720 1277.230 840.000 ;
        RECT 1278.070 835.720 1280.910 840.000 ;
        RECT 1281.750 835.720 1285.050 840.000 ;
        RECT 1285.890 835.720 1288.730 840.000 ;
        RECT 1289.570 835.720 1292.410 840.000 ;
        RECT 1293.250 835.720 1296.090 840.000 ;
        RECT 1296.930 835.720 1299.770 840.000 ;
        RECT 1300.610 835.720 1303.910 840.000 ;
        RECT 1304.750 835.720 1307.590 840.000 ;
        RECT 1308.430 835.720 1311.270 840.000 ;
        RECT 1312.110 835.720 1314.950 840.000 ;
        RECT 1315.790 835.720 1319.090 840.000 ;
        RECT 1319.930 835.720 1322.770 840.000 ;
        RECT 1323.610 835.720 1326.450 840.000 ;
        RECT 1327.290 835.720 1330.130 840.000 ;
        RECT 1330.970 835.720 1333.810 840.000 ;
        RECT 1334.650 835.720 1337.950 840.000 ;
        RECT 1338.790 835.720 1341.630 840.000 ;
        RECT 1342.470 835.720 1345.310 840.000 ;
        RECT 1346.150 835.720 1348.990 840.000 ;
        RECT 1349.830 835.720 1352.670 840.000 ;
        RECT 1353.510 835.720 1356.810 840.000 ;
        RECT 1357.650 835.720 1360.490 840.000 ;
        RECT 1361.330 835.720 1364.170 840.000 ;
        RECT 1365.010 835.720 1367.850 840.000 ;
        RECT 1368.690 835.720 1371.530 840.000 ;
        RECT 1372.370 835.720 1375.670 840.000 ;
        RECT 1376.510 835.720 1379.350 840.000 ;
        RECT 1380.190 835.720 1383.030 840.000 ;
        RECT 1383.870 835.720 1386.710 840.000 ;
        RECT 1387.550 835.720 1390.390 840.000 ;
        RECT 1391.230 835.720 1394.530 840.000 ;
        RECT 1395.370 835.720 1398.210 840.000 ;
        RECT 1399.050 835.720 1401.890 840.000 ;
        RECT 1402.730 835.720 1405.570 840.000 ;
        RECT 1406.410 835.720 1409.250 840.000 ;
        RECT 1410.090 835.720 1413.390 840.000 ;
        RECT 1414.230 835.720 1417.070 840.000 ;
        RECT 1417.910 835.720 1420.750 840.000 ;
        RECT 1421.590 835.720 1424.430 840.000 ;
        RECT 1425.270 835.720 1428.570 840.000 ;
        RECT 1429.410 835.720 1432.250 840.000 ;
        RECT 1433.090 835.720 1435.930 840.000 ;
        RECT 1436.770 835.720 1439.610 840.000 ;
        RECT 1440.450 835.720 1443.290 840.000 ;
        RECT 1444.130 835.720 1447.430 840.000 ;
        RECT 1448.270 835.720 1451.110 840.000 ;
        RECT 1451.950 835.720 1454.790 840.000 ;
        RECT 1455.630 835.720 1458.470 840.000 ;
        RECT 1459.310 835.720 1462.150 840.000 ;
        RECT 1462.990 835.720 1466.290 840.000 ;
        RECT 1467.130 835.720 1469.970 840.000 ;
        RECT 1470.810 835.720 1473.650 840.000 ;
        RECT 1474.490 835.720 1477.330 840.000 ;
        RECT 1478.170 835.720 1481.010 840.000 ;
        RECT 1481.850 835.720 1485.150 840.000 ;
        RECT 1485.990 835.720 1488.830 840.000 ;
        RECT 1489.670 835.720 1492.510 840.000 ;
        RECT 1493.350 835.720 1496.190 840.000 ;
        RECT 1497.030 835.720 1499.870 840.000 ;
        RECT 1500.710 835.720 1504.010 840.000 ;
        RECT 1504.850 835.720 1507.690 840.000 ;
        RECT 1508.530 835.720 1511.370 840.000 ;
        RECT 1512.210 835.720 1515.050 840.000 ;
        RECT 1515.890 835.720 1518.730 840.000 ;
        RECT 1519.570 835.720 1522.870 840.000 ;
        RECT 1523.710 835.720 1526.550 840.000 ;
        RECT 1527.390 835.720 1530.230 840.000 ;
        RECT 1531.070 835.720 1533.910 840.000 ;
        RECT 1534.750 835.720 1537.590 840.000 ;
        RECT 1538.430 835.720 1541.730 840.000 ;
        RECT 1542.570 835.720 1545.410 840.000 ;
        RECT 1546.250 835.720 1549.090 840.000 ;
        RECT 1549.930 835.720 1552.770 840.000 ;
        RECT 1553.610 835.720 1556.910 840.000 ;
        RECT 1557.750 835.720 1560.590 840.000 ;
        RECT 1561.430 835.720 1564.270 840.000 ;
        RECT 1565.110 835.720 1567.950 840.000 ;
        RECT 1568.790 835.720 1571.630 840.000 ;
        RECT 1572.470 835.720 1575.770 840.000 ;
        RECT 1576.610 835.720 1579.450 840.000 ;
        RECT 1580.290 835.720 1583.130 840.000 ;
        RECT 1583.970 835.720 1586.810 840.000 ;
        RECT 1587.650 835.720 1590.490 840.000 ;
        RECT 1591.330 835.720 1594.630 840.000 ;
        RECT 1595.470 835.720 1598.310 840.000 ;
        RECT 1599.150 835.720 1601.990 840.000 ;
        RECT 1602.830 835.720 1605.670 840.000 ;
        RECT 1606.510 835.720 1609.350 840.000 ;
        RECT 1610.190 835.720 1613.490 840.000 ;
        RECT 1614.330 835.720 1617.170 840.000 ;
        RECT 1618.010 835.720 1620.850 840.000 ;
        RECT 1621.690 835.720 1624.530 840.000 ;
        RECT 1625.370 835.720 1628.210 840.000 ;
        RECT 1629.050 835.720 1632.350 840.000 ;
        RECT 1633.190 835.720 1636.030 840.000 ;
        RECT 1636.870 835.720 1639.710 840.000 ;
        RECT 1640.550 835.720 1643.390 840.000 ;
        RECT 1644.230 835.720 1647.070 840.000 ;
        RECT 1647.910 835.720 1651.210 840.000 ;
        RECT 1652.050 835.720 1654.890 840.000 ;
        RECT 1655.730 835.720 1658.570 840.000 ;
        RECT 1659.410 835.720 1662.250 840.000 ;
        RECT 1663.090 835.720 1666.390 840.000 ;
        RECT 1667.230 835.720 1670.070 840.000 ;
        RECT 1670.910 835.720 1673.750 840.000 ;
        RECT 1674.590 835.720 1677.430 840.000 ;
        RECT 1678.270 835.720 1681.110 840.000 ;
        RECT 1681.950 835.720 1685.250 840.000 ;
        RECT 1686.090 835.720 1688.930 840.000 ;
        RECT 1689.770 835.720 1692.610 840.000 ;
        RECT 1693.450 835.720 1696.290 840.000 ;
        RECT 1697.130 835.720 1699.970 840.000 ;
        RECT 1700.810 835.720 1704.110 840.000 ;
        RECT 1704.950 835.720 1707.790 840.000 ;
        RECT 1708.630 835.720 1711.470 840.000 ;
        RECT 1712.310 835.720 1715.150 840.000 ;
        RECT 1715.990 835.720 1718.830 840.000 ;
        RECT 1719.670 835.720 1722.970 840.000 ;
        RECT 1723.810 835.720 1726.650 840.000 ;
        RECT 1727.490 835.720 1730.330 840.000 ;
        RECT 1731.170 835.720 1734.010 840.000 ;
        RECT 1734.850 835.720 1737.690 840.000 ;
        RECT 1738.530 835.720 1741.830 840.000 ;
        RECT 1742.670 835.720 1745.510 840.000 ;
        RECT 1746.350 835.720 1749.190 840.000 ;
        RECT 1750.030 835.720 1752.870 840.000 ;
        RECT 1753.710 835.720 1756.550 840.000 ;
        RECT 1757.390 835.720 1760.690 840.000 ;
        RECT 1761.530 835.720 1764.370 840.000 ;
        RECT 1765.210 835.720 1768.050 840.000 ;
        RECT 1768.890 835.720 1771.730 840.000 ;
        RECT 1772.570 835.720 1775.410 840.000 ;
        RECT 1776.250 835.720 1779.550 840.000 ;
        RECT 1780.390 835.720 1783.230 840.000 ;
        RECT 1784.070 835.720 1786.910 840.000 ;
        RECT 1787.750 835.720 1790.590 840.000 ;
        RECT 1791.430 835.720 1794.730 840.000 ;
        RECT 1795.570 835.720 1798.410 840.000 ;
        RECT 1799.250 835.720 1802.090 840.000 ;
        RECT 1802.930 835.720 1805.770 840.000 ;
        RECT 1806.610 835.720 1809.450 840.000 ;
        RECT 1810.290 835.720 1813.590 840.000 ;
        RECT 1814.430 835.720 1817.270 840.000 ;
        RECT 1818.110 835.720 1820.950 840.000 ;
        RECT 1821.790 835.720 1824.630 840.000 ;
        RECT 1825.470 835.720 1828.310 840.000 ;
        RECT 1829.150 835.720 1832.450 840.000 ;
        RECT 1833.290 835.720 1836.130 840.000 ;
        RECT 1836.970 835.720 1839.810 840.000 ;
        RECT 1840.650 835.720 1843.490 840.000 ;
        RECT 1844.330 835.720 1847.170 840.000 ;
        RECT 1848.010 835.720 1851.310 840.000 ;
        RECT 1852.150 835.720 1854.990 840.000 ;
        RECT 1855.830 835.720 1858.670 840.000 ;
        RECT 1859.510 835.720 1862.350 840.000 ;
        RECT 1863.190 835.720 1866.030 840.000 ;
        RECT 1866.870 835.720 1870.170 840.000 ;
        RECT 1871.010 835.720 1873.850 840.000 ;
        RECT 1874.690 835.720 1877.530 840.000 ;
        RECT 1878.370 835.720 1881.210 840.000 ;
        RECT 1882.050 835.720 1884.890 840.000 ;
        RECT 1885.730 835.720 1889.030 840.000 ;
        RECT 1889.870 835.720 1892.710 840.000 ;
        RECT 1893.550 835.720 1896.390 840.000 ;
        RECT 1897.230 835.720 1900.070 840.000 ;
        RECT 1900.910 835.720 1904.210 840.000 ;
        RECT 1905.050 835.720 1907.890 840.000 ;
        RECT 1908.730 835.720 1911.570 840.000 ;
        RECT 1912.410 835.720 1915.250 840.000 ;
        RECT 1916.090 835.720 1918.930 840.000 ;
        RECT 1919.770 835.720 1923.070 840.000 ;
        RECT 1923.910 835.720 1926.750 840.000 ;
        RECT 1927.590 835.720 1930.430 840.000 ;
        RECT 1931.270 835.720 1934.110 840.000 ;
        RECT 1934.950 835.720 1937.790 840.000 ;
        RECT 1938.630 835.720 1941.930 840.000 ;
        RECT 1942.770 835.720 1945.610 840.000 ;
        RECT 1946.450 835.720 1949.290 840.000 ;
        RECT 1950.130 835.720 1952.970 840.000 ;
        RECT 1953.810 835.720 1956.650 840.000 ;
        RECT 1957.490 835.720 1960.790 840.000 ;
        RECT 1961.630 835.720 1964.470 840.000 ;
        RECT 1965.310 835.720 1968.150 840.000 ;
        RECT 1968.990 835.720 1971.830 840.000 ;
        RECT 1972.670 835.720 1975.510 840.000 ;
        RECT 1976.350 835.720 1979.650 840.000 ;
        RECT 1980.490 835.720 1983.330 840.000 ;
        RECT 1984.170 835.720 1987.010 840.000 ;
        RECT 1987.850 835.720 1990.690 840.000 ;
        RECT 1991.530 835.720 1994.370 840.000 ;
        RECT 1995.210 835.720 1998.510 840.000 ;
        RECT 1999.350 835.720 2002.190 840.000 ;
        RECT 2003.030 835.720 2005.870 840.000 ;
        RECT 2006.710 835.720 2009.550 840.000 ;
        RECT 2010.390 835.720 2013.230 840.000 ;
        RECT 2014.070 835.720 2017.370 840.000 ;
        RECT 2018.210 835.720 2021.050 840.000 ;
        RECT 2021.890 835.720 2024.730 840.000 ;
        RECT 2025.570 835.720 2028.410 840.000 ;
        RECT 2029.250 835.720 2032.550 840.000 ;
        RECT 2033.390 835.720 2036.230 840.000 ;
        RECT 2037.070 835.720 2039.910 840.000 ;
        RECT 2040.750 835.720 2043.590 840.000 ;
        RECT 2044.430 835.720 2047.270 840.000 ;
        RECT 2048.110 835.720 2051.410 840.000 ;
        RECT 2052.250 835.720 2055.090 840.000 ;
        RECT 2055.930 835.720 2058.770 840.000 ;
        RECT 2059.610 835.720 2062.450 840.000 ;
        RECT 2063.290 835.720 2066.130 840.000 ;
        RECT 2066.970 835.720 2070.270 840.000 ;
        RECT 2071.110 835.720 2073.950 840.000 ;
        RECT 2074.790 835.720 2077.630 840.000 ;
        RECT 2078.470 835.720 2081.310 840.000 ;
        RECT 2082.150 835.720 2084.990 840.000 ;
        RECT 2085.830 835.720 2089.130 840.000 ;
        RECT 2089.970 835.720 2092.810 840.000 ;
        RECT 2093.650 835.720 2096.490 840.000 ;
        RECT 2097.330 835.720 2100.170 840.000 ;
        RECT 2101.010 835.720 2103.850 840.000 ;
        RECT 2104.690 835.720 2107.990 840.000 ;
        RECT 2108.830 835.720 2111.670 840.000 ;
        RECT 2112.510 835.720 2115.350 840.000 ;
        RECT 2116.190 835.720 2119.030 840.000 ;
        RECT 2119.870 835.720 2122.710 840.000 ;
        RECT 2123.550 835.720 2126.850 840.000 ;
        RECT 2127.690 835.720 2130.530 840.000 ;
        RECT 2131.370 835.720 2134.210 840.000 ;
        RECT 2135.050 835.720 2137.890 840.000 ;
        RECT 2138.730 835.720 2142.030 840.000 ;
        RECT 2142.870 835.720 2145.710 840.000 ;
        RECT 2146.550 835.720 2149.390 840.000 ;
        RECT 2150.230 835.720 2153.070 840.000 ;
        RECT 2153.910 835.720 2156.750 840.000 ;
        RECT 2157.590 835.720 2160.890 840.000 ;
        RECT 2161.730 835.720 2164.570 840.000 ;
        RECT 2165.410 835.720 2168.250 840.000 ;
        RECT 2169.090 835.720 2171.930 840.000 ;
        RECT 2172.770 835.720 2175.610 840.000 ;
        RECT 2176.450 835.720 2179.750 840.000 ;
        RECT 2180.590 835.720 2183.430 840.000 ;
        RECT 2184.270 835.720 2187.110 840.000 ;
        RECT 2187.950 835.720 2190.790 840.000 ;
        RECT 2191.630 835.720 2194.470 840.000 ;
        RECT 2195.310 835.720 2198.610 840.000 ;
        RECT 2199.450 835.720 2202.290 840.000 ;
        RECT 2203.130 835.720 2205.970 840.000 ;
        RECT 2206.810 835.720 2209.650 840.000 ;
        RECT 2210.490 835.720 2213.330 840.000 ;
        RECT 2214.170 835.720 2217.470 840.000 ;
        RECT 2218.310 835.720 2221.150 840.000 ;
        RECT 2221.990 835.720 2224.830 840.000 ;
        RECT 2225.670 835.720 2228.510 840.000 ;
        RECT 2229.350 835.720 2232.190 840.000 ;
        RECT 2233.030 835.720 2236.330 840.000 ;
        RECT 2237.170 835.720 2240.010 840.000 ;
        RECT 2240.850 835.720 2243.690 840.000 ;
        RECT 2244.530 835.720 2247.370 840.000 ;
        RECT 0.090 4.280 2247.860 835.720 ;
        RECT 0.090 4.000 43.050 4.280 ;
        RECT 43.890 4.000 129.530 4.280 ;
        RECT 130.370 4.000 216.010 4.280 ;
        RECT 216.850 4.000 302.490 4.280 ;
        RECT 303.330 4.000 388.970 4.280 ;
        RECT 389.810 4.000 475.450 4.280 ;
        RECT 476.290 4.000 561.930 4.280 ;
        RECT 562.770 4.000 648.410 4.280 ;
        RECT 649.250 4.000 734.890 4.280 ;
        RECT 735.730 4.000 821.830 4.280 ;
        RECT 822.670 4.000 908.310 4.280 ;
        RECT 909.150 4.000 994.790 4.280 ;
        RECT 995.630 4.000 1081.270 4.280 ;
        RECT 1082.110 4.000 1167.750 4.280 ;
        RECT 1168.590 4.000 1254.230 4.280 ;
        RECT 1255.070 4.000 1340.710 4.280 ;
        RECT 1341.550 4.000 1427.190 4.280 ;
        RECT 1428.030 4.000 1513.670 4.280 ;
        RECT 1514.510 4.000 1600.610 4.280 ;
        RECT 1601.450 4.000 1687.090 4.280 ;
        RECT 1687.930 4.000 1773.570 4.280 ;
        RECT 1774.410 4.000 1860.050 4.280 ;
        RECT 1860.890 4.000 1946.530 4.280 ;
        RECT 1947.370 4.000 2033.010 4.280 ;
        RECT 2033.850 4.000 2119.490 4.280 ;
        RECT 2120.330 4.000 2205.970 4.280 ;
        RECT 2206.810 4.000 2247.860 4.280 ;
      LAYER met3 ;
        RECT 4.400 836.720 2246.000 837.585 ;
        RECT 0.065 835.400 2246.000 836.720 ;
        RECT 0.065 834.040 2245.600 835.400 ;
        RECT 4.400 834.000 2245.600 834.040 ;
        RECT 4.400 832.640 2246.000 834.000 ;
        RECT 0.065 830.640 2246.000 832.640 ;
        RECT 4.400 829.240 2246.000 830.640 ;
        RECT 0.065 826.560 2246.000 829.240 ;
        RECT 4.400 825.880 2246.000 826.560 ;
        RECT 4.400 825.160 2245.600 825.880 ;
        RECT 0.065 824.480 2245.600 825.160 ;
        RECT 0.065 823.160 2246.000 824.480 ;
        RECT 4.400 821.760 2246.000 823.160 ;
        RECT 0.065 819.080 2246.000 821.760 ;
        RECT 4.400 817.680 2246.000 819.080 ;
        RECT 0.065 816.360 2246.000 817.680 ;
        RECT 0.065 815.000 2245.600 816.360 ;
        RECT 4.400 814.960 2245.600 815.000 ;
        RECT 4.400 813.600 2246.000 814.960 ;
        RECT 0.065 811.600 2246.000 813.600 ;
        RECT 4.400 810.200 2246.000 811.600 ;
        RECT 0.065 807.520 2246.000 810.200 ;
        RECT 4.400 806.840 2246.000 807.520 ;
        RECT 4.400 806.120 2245.600 806.840 ;
        RECT 0.065 805.440 2245.600 806.120 ;
        RECT 0.065 804.120 2246.000 805.440 ;
        RECT 4.400 802.720 2246.000 804.120 ;
        RECT 0.065 800.040 2246.000 802.720 ;
        RECT 4.400 798.640 2246.000 800.040 ;
        RECT 0.065 797.320 2246.000 798.640 ;
        RECT 0.065 795.960 2245.600 797.320 ;
        RECT 4.400 795.920 2245.600 795.960 ;
        RECT 4.400 794.560 2246.000 795.920 ;
        RECT 0.065 792.560 2246.000 794.560 ;
        RECT 4.400 791.160 2246.000 792.560 ;
        RECT 0.065 788.480 2246.000 791.160 ;
        RECT 4.400 787.800 2246.000 788.480 ;
        RECT 4.400 787.080 2245.600 787.800 ;
        RECT 0.065 786.400 2245.600 787.080 ;
        RECT 0.065 785.080 2246.000 786.400 ;
        RECT 4.400 783.680 2246.000 785.080 ;
        RECT 0.065 781.000 2246.000 783.680 ;
        RECT 4.400 779.600 2246.000 781.000 ;
        RECT 0.065 778.280 2246.000 779.600 ;
        RECT 0.065 777.600 2245.600 778.280 ;
        RECT 4.400 776.880 2245.600 777.600 ;
        RECT 4.400 776.200 2246.000 776.880 ;
        RECT 0.065 773.520 2246.000 776.200 ;
        RECT 4.400 772.120 2246.000 773.520 ;
        RECT 0.065 769.440 2246.000 772.120 ;
        RECT 4.400 768.760 2246.000 769.440 ;
        RECT 4.400 768.040 2245.600 768.760 ;
        RECT 0.065 767.360 2245.600 768.040 ;
        RECT 0.065 766.040 2246.000 767.360 ;
        RECT 4.400 764.640 2246.000 766.040 ;
        RECT 0.065 761.960 2246.000 764.640 ;
        RECT 4.400 760.560 2246.000 761.960 ;
        RECT 0.065 759.240 2246.000 760.560 ;
        RECT 0.065 758.560 2245.600 759.240 ;
        RECT 4.400 757.840 2245.600 758.560 ;
        RECT 4.400 757.160 2246.000 757.840 ;
        RECT 0.065 754.480 2246.000 757.160 ;
        RECT 4.400 753.080 2246.000 754.480 ;
        RECT 0.065 750.400 2246.000 753.080 ;
        RECT 4.400 749.720 2246.000 750.400 ;
        RECT 4.400 749.000 2245.600 749.720 ;
        RECT 0.065 748.320 2245.600 749.000 ;
        RECT 0.065 747.000 2246.000 748.320 ;
        RECT 4.400 745.600 2246.000 747.000 ;
        RECT 0.065 742.920 2246.000 745.600 ;
        RECT 4.400 741.520 2246.000 742.920 ;
        RECT 0.065 740.200 2246.000 741.520 ;
        RECT 0.065 739.520 2245.600 740.200 ;
        RECT 4.400 738.800 2245.600 739.520 ;
        RECT 4.400 738.120 2246.000 738.800 ;
        RECT 0.065 735.440 2246.000 738.120 ;
        RECT 4.400 734.040 2246.000 735.440 ;
        RECT 0.065 731.360 2246.000 734.040 ;
        RECT 4.400 730.680 2246.000 731.360 ;
        RECT 4.400 729.960 2245.600 730.680 ;
        RECT 0.065 729.280 2245.600 729.960 ;
        RECT 0.065 727.960 2246.000 729.280 ;
        RECT 4.400 726.560 2246.000 727.960 ;
        RECT 0.065 723.880 2246.000 726.560 ;
        RECT 4.400 722.480 2246.000 723.880 ;
        RECT 0.065 721.160 2246.000 722.480 ;
        RECT 0.065 720.480 2245.600 721.160 ;
        RECT 4.400 719.760 2245.600 720.480 ;
        RECT 4.400 719.080 2246.000 719.760 ;
        RECT 0.065 716.400 2246.000 719.080 ;
        RECT 4.400 715.000 2246.000 716.400 ;
        RECT 0.065 713.000 2246.000 715.000 ;
        RECT 4.400 711.640 2246.000 713.000 ;
        RECT 4.400 711.600 2245.600 711.640 ;
        RECT 0.065 710.240 2245.600 711.600 ;
        RECT 0.065 708.920 2246.000 710.240 ;
        RECT 4.400 707.520 2246.000 708.920 ;
        RECT 0.065 704.840 2246.000 707.520 ;
        RECT 4.400 703.440 2246.000 704.840 ;
        RECT 0.065 702.120 2246.000 703.440 ;
        RECT 0.065 701.440 2245.600 702.120 ;
        RECT 4.400 700.720 2245.600 701.440 ;
        RECT 4.400 700.040 2246.000 700.720 ;
        RECT 0.065 697.360 2246.000 700.040 ;
        RECT 4.400 695.960 2246.000 697.360 ;
        RECT 0.065 693.960 2246.000 695.960 ;
        RECT 4.400 692.600 2246.000 693.960 ;
        RECT 4.400 692.560 2245.600 692.600 ;
        RECT 0.065 691.200 2245.600 692.560 ;
        RECT 0.065 689.880 2246.000 691.200 ;
        RECT 4.400 688.480 2246.000 689.880 ;
        RECT 0.065 685.800 2246.000 688.480 ;
        RECT 4.400 684.400 2246.000 685.800 ;
        RECT 0.065 683.080 2246.000 684.400 ;
        RECT 0.065 682.400 2245.600 683.080 ;
        RECT 4.400 681.680 2245.600 682.400 ;
        RECT 4.400 681.000 2246.000 681.680 ;
        RECT 0.065 678.320 2246.000 681.000 ;
        RECT 4.400 676.920 2246.000 678.320 ;
        RECT 0.065 674.920 2246.000 676.920 ;
        RECT 4.400 673.560 2246.000 674.920 ;
        RECT 4.400 673.520 2245.600 673.560 ;
        RECT 0.065 672.160 2245.600 673.520 ;
        RECT 0.065 670.840 2246.000 672.160 ;
        RECT 4.400 669.440 2246.000 670.840 ;
        RECT 0.065 666.760 2246.000 669.440 ;
        RECT 4.400 665.360 2246.000 666.760 ;
        RECT 0.065 664.040 2246.000 665.360 ;
        RECT 0.065 663.360 2245.600 664.040 ;
        RECT 4.400 662.640 2245.600 663.360 ;
        RECT 4.400 661.960 2246.000 662.640 ;
        RECT 0.065 659.280 2246.000 661.960 ;
        RECT 4.400 657.880 2246.000 659.280 ;
        RECT 0.065 655.880 2246.000 657.880 ;
        RECT 4.400 654.520 2246.000 655.880 ;
        RECT 4.400 654.480 2245.600 654.520 ;
        RECT 0.065 653.120 2245.600 654.480 ;
        RECT 0.065 651.800 2246.000 653.120 ;
        RECT 4.400 650.400 2246.000 651.800 ;
        RECT 0.065 648.400 2246.000 650.400 ;
        RECT 4.400 647.000 2246.000 648.400 ;
        RECT 0.065 645.000 2246.000 647.000 ;
        RECT 0.065 644.320 2245.600 645.000 ;
        RECT 4.400 643.600 2245.600 644.320 ;
        RECT 4.400 642.920 2246.000 643.600 ;
        RECT 0.065 640.240 2246.000 642.920 ;
        RECT 4.400 638.840 2246.000 640.240 ;
        RECT 0.065 636.840 2246.000 638.840 ;
        RECT 4.400 635.480 2246.000 636.840 ;
        RECT 4.400 635.440 2245.600 635.480 ;
        RECT 0.065 634.080 2245.600 635.440 ;
        RECT 0.065 632.760 2246.000 634.080 ;
        RECT 4.400 631.360 2246.000 632.760 ;
        RECT 0.065 629.360 2246.000 631.360 ;
        RECT 4.400 627.960 2246.000 629.360 ;
        RECT 0.065 625.960 2246.000 627.960 ;
        RECT 0.065 625.280 2245.600 625.960 ;
        RECT 4.400 624.560 2245.600 625.280 ;
        RECT 4.400 623.880 2246.000 624.560 ;
        RECT 0.065 621.200 2246.000 623.880 ;
        RECT 4.400 619.800 2246.000 621.200 ;
        RECT 0.065 617.800 2246.000 619.800 ;
        RECT 4.400 616.440 2246.000 617.800 ;
        RECT 4.400 616.400 2245.600 616.440 ;
        RECT 0.065 615.040 2245.600 616.400 ;
        RECT 0.065 613.720 2246.000 615.040 ;
        RECT 4.400 612.320 2246.000 613.720 ;
        RECT 0.065 610.320 2246.000 612.320 ;
        RECT 4.400 608.920 2246.000 610.320 ;
        RECT 0.065 606.920 2246.000 608.920 ;
        RECT 0.065 606.240 2245.600 606.920 ;
        RECT 4.400 605.520 2245.600 606.240 ;
        RECT 4.400 604.840 2246.000 605.520 ;
        RECT 0.065 602.160 2246.000 604.840 ;
        RECT 4.400 600.760 2246.000 602.160 ;
        RECT 0.065 598.760 2246.000 600.760 ;
        RECT 4.400 597.400 2246.000 598.760 ;
        RECT 4.400 597.360 2245.600 597.400 ;
        RECT 0.065 596.000 2245.600 597.360 ;
        RECT 0.065 594.680 2246.000 596.000 ;
        RECT 4.400 593.280 2246.000 594.680 ;
        RECT 0.065 591.280 2246.000 593.280 ;
        RECT 4.400 589.880 2246.000 591.280 ;
        RECT 0.065 587.880 2246.000 589.880 ;
        RECT 0.065 587.200 2245.600 587.880 ;
        RECT 4.400 586.480 2245.600 587.200 ;
        RECT 4.400 585.800 2246.000 586.480 ;
        RECT 0.065 583.800 2246.000 585.800 ;
        RECT 4.400 582.400 2246.000 583.800 ;
        RECT 0.065 579.720 2246.000 582.400 ;
        RECT 4.400 578.360 2246.000 579.720 ;
        RECT 4.400 578.320 2245.600 578.360 ;
        RECT 0.065 576.960 2245.600 578.320 ;
        RECT 0.065 575.640 2246.000 576.960 ;
        RECT 4.400 574.240 2246.000 575.640 ;
        RECT 0.065 572.240 2246.000 574.240 ;
        RECT 4.400 570.840 2246.000 572.240 ;
        RECT 0.065 568.840 2246.000 570.840 ;
        RECT 0.065 568.160 2245.600 568.840 ;
        RECT 4.400 567.440 2245.600 568.160 ;
        RECT 4.400 566.760 2246.000 567.440 ;
        RECT 0.065 564.760 2246.000 566.760 ;
        RECT 4.400 563.360 2246.000 564.760 ;
        RECT 0.065 560.680 2246.000 563.360 ;
        RECT 4.400 559.280 2246.000 560.680 ;
        RECT 0.065 558.640 2246.000 559.280 ;
        RECT 0.065 557.240 2245.600 558.640 ;
        RECT 0.065 556.600 2246.000 557.240 ;
        RECT 4.400 555.200 2246.000 556.600 ;
        RECT 0.065 553.200 2246.000 555.200 ;
        RECT 4.400 551.800 2246.000 553.200 ;
        RECT 0.065 549.120 2246.000 551.800 ;
        RECT 4.400 547.720 2245.600 549.120 ;
        RECT 0.065 545.720 2246.000 547.720 ;
        RECT 4.400 544.320 2246.000 545.720 ;
        RECT 0.065 541.640 2246.000 544.320 ;
        RECT 4.400 540.240 2246.000 541.640 ;
        RECT 0.065 539.600 2246.000 540.240 ;
        RECT 0.065 538.200 2245.600 539.600 ;
        RECT 0.065 537.560 2246.000 538.200 ;
        RECT 4.400 536.160 2246.000 537.560 ;
        RECT 0.065 534.160 2246.000 536.160 ;
        RECT 4.400 532.760 2246.000 534.160 ;
        RECT 0.065 530.080 2246.000 532.760 ;
        RECT 4.400 528.680 2245.600 530.080 ;
        RECT 0.065 526.680 2246.000 528.680 ;
        RECT 4.400 525.280 2246.000 526.680 ;
        RECT 0.065 522.600 2246.000 525.280 ;
        RECT 4.400 521.200 2246.000 522.600 ;
        RECT 0.065 520.560 2246.000 521.200 ;
        RECT 0.065 519.200 2245.600 520.560 ;
        RECT 4.400 519.160 2245.600 519.200 ;
        RECT 4.400 517.800 2246.000 519.160 ;
        RECT 0.065 515.120 2246.000 517.800 ;
        RECT 4.400 513.720 2246.000 515.120 ;
        RECT 0.065 511.040 2246.000 513.720 ;
        RECT 4.400 509.640 2245.600 511.040 ;
        RECT 0.065 507.640 2246.000 509.640 ;
        RECT 4.400 506.240 2246.000 507.640 ;
        RECT 0.065 503.560 2246.000 506.240 ;
        RECT 4.400 502.160 2246.000 503.560 ;
        RECT 0.065 501.520 2246.000 502.160 ;
        RECT 0.065 500.160 2245.600 501.520 ;
        RECT 4.400 500.120 2245.600 500.160 ;
        RECT 4.400 498.760 2246.000 500.120 ;
        RECT 0.065 496.080 2246.000 498.760 ;
        RECT 4.400 494.680 2246.000 496.080 ;
        RECT 0.065 492.000 2246.000 494.680 ;
        RECT 4.400 490.600 2245.600 492.000 ;
        RECT 0.065 488.600 2246.000 490.600 ;
        RECT 4.400 487.200 2246.000 488.600 ;
        RECT 0.065 484.520 2246.000 487.200 ;
        RECT 4.400 483.120 2246.000 484.520 ;
        RECT 0.065 482.480 2246.000 483.120 ;
        RECT 0.065 481.120 2245.600 482.480 ;
        RECT 4.400 481.080 2245.600 481.120 ;
        RECT 4.400 479.720 2246.000 481.080 ;
        RECT 0.065 477.040 2246.000 479.720 ;
        RECT 4.400 475.640 2246.000 477.040 ;
        RECT 0.065 472.960 2246.000 475.640 ;
        RECT 4.400 471.560 2245.600 472.960 ;
        RECT 0.065 469.560 2246.000 471.560 ;
        RECT 4.400 468.160 2246.000 469.560 ;
        RECT 0.065 465.480 2246.000 468.160 ;
        RECT 4.400 464.080 2246.000 465.480 ;
        RECT 0.065 463.440 2246.000 464.080 ;
        RECT 0.065 462.080 2245.600 463.440 ;
        RECT 4.400 462.040 2245.600 462.080 ;
        RECT 4.400 460.680 2246.000 462.040 ;
        RECT 0.065 458.000 2246.000 460.680 ;
        RECT 4.400 456.600 2246.000 458.000 ;
        RECT 0.065 454.600 2246.000 456.600 ;
        RECT 4.400 453.920 2246.000 454.600 ;
        RECT 4.400 453.200 2245.600 453.920 ;
        RECT 0.065 452.520 2245.600 453.200 ;
        RECT 0.065 450.520 2246.000 452.520 ;
        RECT 4.400 449.120 2246.000 450.520 ;
        RECT 0.065 446.440 2246.000 449.120 ;
        RECT 4.400 445.040 2246.000 446.440 ;
        RECT 0.065 444.400 2246.000 445.040 ;
        RECT 0.065 443.040 2245.600 444.400 ;
        RECT 4.400 443.000 2245.600 443.040 ;
        RECT 4.400 441.640 2246.000 443.000 ;
        RECT 0.065 438.960 2246.000 441.640 ;
        RECT 4.400 437.560 2246.000 438.960 ;
        RECT 0.065 435.560 2246.000 437.560 ;
        RECT 4.400 434.880 2246.000 435.560 ;
        RECT 4.400 434.160 2245.600 434.880 ;
        RECT 0.065 433.480 2245.600 434.160 ;
        RECT 0.065 431.480 2246.000 433.480 ;
        RECT 4.400 430.080 2246.000 431.480 ;
        RECT 0.065 427.400 2246.000 430.080 ;
        RECT 4.400 426.000 2246.000 427.400 ;
        RECT 0.065 425.360 2246.000 426.000 ;
        RECT 0.065 424.000 2245.600 425.360 ;
        RECT 4.400 423.960 2245.600 424.000 ;
        RECT 4.400 422.600 2246.000 423.960 ;
        RECT 0.065 419.920 2246.000 422.600 ;
        RECT 4.400 418.520 2246.000 419.920 ;
        RECT 0.065 416.520 2246.000 418.520 ;
        RECT 4.400 415.840 2246.000 416.520 ;
        RECT 4.400 415.120 2245.600 415.840 ;
        RECT 0.065 414.440 2245.600 415.120 ;
        RECT 0.065 412.440 2246.000 414.440 ;
        RECT 4.400 411.040 2246.000 412.440 ;
        RECT 0.065 408.360 2246.000 411.040 ;
        RECT 4.400 406.960 2246.000 408.360 ;
        RECT 0.065 406.320 2246.000 406.960 ;
        RECT 0.065 404.960 2245.600 406.320 ;
        RECT 4.400 404.920 2245.600 404.960 ;
        RECT 4.400 403.560 2246.000 404.920 ;
        RECT 0.065 400.880 2246.000 403.560 ;
        RECT 4.400 399.480 2246.000 400.880 ;
        RECT 0.065 397.480 2246.000 399.480 ;
        RECT 4.400 396.800 2246.000 397.480 ;
        RECT 4.400 396.080 2245.600 396.800 ;
        RECT 0.065 395.400 2245.600 396.080 ;
        RECT 0.065 393.400 2246.000 395.400 ;
        RECT 4.400 392.000 2246.000 393.400 ;
        RECT 0.065 390.000 2246.000 392.000 ;
        RECT 4.400 388.600 2246.000 390.000 ;
        RECT 0.065 387.280 2246.000 388.600 ;
        RECT 0.065 385.920 2245.600 387.280 ;
        RECT 4.400 385.880 2245.600 385.920 ;
        RECT 4.400 384.520 2246.000 385.880 ;
        RECT 0.065 381.840 2246.000 384.520 ;
        RECT 4.400 380.440 2246.000 381.840 ;
        RECT 0.065 378.440 2246.000 380.440 ;
        RECT 4.400 377.760 2246.000 378.440 ;
        RECT 4.400 377.040 2245.600 377.760 ;
        RECT 0.065 376.360 2245.600 377.040 ;
        RECT 0.065 374.360 2246.000 376.360 ;
        RECT 4.400 372.960 2246.000 374.360 ;
        RECT 0.065 370.960 2246.000 372.960 ;
        RECT 4.400 369.560 2246.000 370.960 ;
        RECT 0.065 368.240 2246.000 369.560 ;
        RECT 0.065 366.880 2245.600 368.240 ;
        RECT 4.400 366.840 2245.600 366.880 ;
        RECT 4.400 365.480 2246.000 366.840 ;
        RECT 0.065 362.800 2246.000 365.480 ;
        RECT 4.400 361.400 2246.000 362.800 ;
        RECT 0.065 359.400 2246.000 361.400 ;
        RECT 4.400 358.720 2246.000 359.400 ;
        RECT 4.400 358.000 2245.600 358.720 ;
        RECT 0.065 357.320 2245.600 358.000 ;
        RECT 0.065 355.320 2246.000 357.320 ;
        RECT 4.400 353.920 2246.000 355.320 ;
        RECT 0.065 351.920 2246.000 353.920 ;
        RECT 4.400 350.520 2246.000 351.920 ;
        RECT 0.065 349.200 2246.000 350.520 ;
        RECT 0.065 347.840 2245.600 349.200 ;
        RECT 4.400 347.800 2245.600 347.840 ;
        RECT 4.400 346.440 2246.000 347.800 ;
        RECT 0.065 343.760 2246.000 346.440 ;
        RECT 4.400 342.360 2246.000 343.760 ;
        RECT 0.065 340.360 2246.000 342.360 ;
        RECT 4.400 339.680 2246.000 340.360 ;
        RECT 4.400 338.960 2245.600 339.680 ;
        RECT 0.065 338.280 2245.600 338.960 ;
        RECT 0.065 336.280 2246.000 338.280 ;
        RECT 4.400 334.880 2246.000 336.280 ;
        RECT 0.065 332.880 2246.000 334.880 ;
        RECT 4.400 331.480 2246.000 332.880 ;
        RECT 0.065 330.160 2246.000 331.480 ;
        RECT 0.065 328.800 2245.600 330.160 ;
        RECT 4.400 328.760 2245.600 328.800 ;
        RECT 4.400 327.400 2246.000 328.760 ;
        RECT 0.065 325.400 2246.000 327.400 ;
        RECT 4.400 324.000 2246.000 325.400 ;
        RECT 0.065 321.320 2246.000 324.000 ;
        RECT 4.400 320.640 2246.000 321.320 ;
        RECT 4.400 319.920 2245.600 320.640 ;
        RECT 0.065 319.240 2245.600 319.920 ;
        RECT 0.065 317.240 2246.000 319.240 ;
        RECT 4.400 315.840 2246.000 317.240 ;
        RECT 0.065 313.840 2246.000 315.840 ;
        RECT 4.400 312.440 2246.000 313.840 ;
        RECT 0.065 311.120 2246.000 312.440 ;
        RECT 0.065 309.760 2245.600 311.120 ;
        RECT 4.400 309.720 2245.600 309.760 ;
        RECT 4.400 308.360 2246.000 309.720 ;
        RECT 0.065 306.360 2246.000 308.360 ;
        RECT 4.400 304.960 2246.000 306.360 ;
        RECT 0.065 302.280 2246.000 304.960 ;
        RECT 4.400 301.600 2246.000 302.280 ;
        RECT 4.400 300.880 2245.600 301.600 ;
        RECT 0.065 300.200 2245.600 300.880 ;
        RECT 0.065 298.200 2246.000 300.200 ;
        RECT 4.400 296.800 2246.000 298.200 ;
        RECT 0.065 294.800 2246.000 296.800 ;
        RECT 4.400 293.400 2246.000 294.800 ;
        RECT 0.065 292.080 2246.000 293.400 ;
        RECT 0.065 290.720 2245.600 292.080 ;
        RECT 4.400 290.680 2245.600 290.720 ;
        RECT 4.400 289.320 2246.000 290.680 ;
        RECT 0.065 287.320 2246.000 289.320 ;
        RECT 4.400 285.920 2246.000 287.320 ;
        RECT 0.065 283.240 2246.000 285.920 ;
        RECT 4.400 281.880 2246.000 283.240 ;
        RECT 4.400 281.840 2245.600 281.880 ;
        RECT 0.065 280.480 2245.600 281.840 ;
        RECT 0.065 279.160 2246.000 280.480 ;
        RECT 4.400 277.760 2246.000 279.160 ;
        RECT 0.065 275.760 2246.000 277.760 ;
        RECT 4.400 274.360 2246.000 275.760 ;
        RECT 0.065 272.360 2246.000 274.360 ;
        RECT 0.065 271.680 2245.600 272.360 ;
        RECT 4.400 270.960 2245.600 271.680 ;
        RECT 4.400 270.280 2246.000 270.960 ;
        RECT 0.065 268.280 2246.000 270.280 ;
        RECT 4.400 266.880 2246.000 268.280 ;
        RECT 0.065 264.200 2246.000 266.880 ;
        RECT 4.400 262.840 2246.000 264.200 ;
        RECT 4.400 262.800 2245.600 262.840 ;
        RECT 0.065 261.440 2245.600 262.800 ;
        RECT 0.065 260.800 2246.000 261.440 ;
        RECT 4.400 259.400 2246.000 260.800 ;
        RECT 0.065 256.720 2246.000 259.400 ;
        RECT 4.400 255.320 2246.000 256.720 ;
        RECT 0.065 253.320 2246.000 255.320 ;
        RECT 0.065 252.640 2245.600 253.320 ;
        RECT 4.400 251.920 2245.600 252.640 ;
        RECT 4.400 251.240 2246.000 251.920 ;
        RECT 0.065 249.240 2246.000 251.240 ;
        RECT 4.400 247.840 2246.000 249.240 ;
        RECT 0.065 245.160 2246.000 247.840 ;
        RECT 4.400 243.800 2246.000 245.160 ;
        RECT 4.400 243.760 2245.600 243.800 ;
        RECT 0.065 242.400 2245.600 243.760 ;
        RECT 0.065 241.760 2246.000 242.400 ;
        RECT 4.400 240.360 2246.000 241.760 ;
        RECT 0.065 237.680 2246.000 240.360 ;
        RECT 4.400 236.280 2246.000 237.680 ;
        RECT 0.065 234.280 2246.000 236.280 ;
        RECT 0.065 233.600 2245.600 234.280 ;
        RECT 4.400 232.880 2245.600 233.600 ;
        RECT 4.400 232.200 2246.000 232.880 ;
        RECT 0.065 230.200 2246.000 232.200 ;
        RECT 4.400 228.800 2246.000 230.200 ;
        RECT 0.065 226.120 2246.000 228.800 ;
        RECT 4.400 224.760 2246.000 226.120 ;
        RECT 4.400 224.720 2245.600 224.760 ;
        RECT 0.065 223.360 2245.600 224.720 ;
        RECT 0.065 222.720 2246.000 223.360 ;
        RECT 4.400 221.320 2246.000 222.720 ;
        RECT 0.065 218.640 2246.000 221.320 ;
        RECT 4.400 217.240 2246.000 218.640 ;
        RECT 0.065 215.240 2246.000 217.240 ;
        RECT 0.065 214.560 2245.600 215.240 ;
        RECT 4.400 213.840 2245.600 214.560 ;
        RECT 4.400 213.160 2246.000 213.840 ;
        RECT 0.065 211.160 2246.000 213.160 ;
        RECT 4.400 209.760 2246.000 211.160 ;
        RECT 0.065 207.080 2246.000 209.760 ;
        RECT 4.400 205.720 2246.000 207.080 ;
        RECT 4.400 205.680 2245.600 205.720 ;
        RECT 0.065 204.320 2245.600 205.680 ;
        RECT 0.065 203.680 2246.000 204.320 ;
        RECT 4.400 202.280 2246.000 203.680 ;
        RECT 0.065 199.600 2246.000 202.280 ;
        RECT 4.400 198.200 2246.000 199.600 ;
        RECT 0.065 196.200 2246.000 198.200 ;
        RECT 4.400 194.800 2245.600 196.200 ;
        RECT 0.065 192.120 2246.000 194.800 ;
        RECT 4.400 190.720 2246.000 192.120 ;
        RECT 0.065 188.040 2246.000 190.720 ;
        RECT 4.400 186.680 2246.000 188.040 ;
        RECT 4.400 186.640 2245.600 186.680 ;
        RECT 0.065 185.280 2245.600 186.640 ;
        RECT 0.065 184.640 2246.000 185.280 ;
        RECT 4.400 183.240 2246.000 184.640 ;
        RECT 0.065 180.560 2246.000 183.240 ;
        RECT 4.400 179.160 2246.000 180.560 ;
        RECT 0.065 177.160 2246.000 179.160 ;
        RECT 4.400 175.760 2245.600 177.160 ;
        RECT 0.065 173.080 2246.000 175.760 ;
        RECT 4.400 171.680 2246.000 173.080 ;
        RECT 0.065 169.000 2246.000 171.680 ;
        RECT 4.400 167.640 2246.000 169.000 ;
        RECT 4.400 167.600 2245.600 167.640 ;
        RECT 0.065 166.240 2245.600 167.600 ;
        RECT 0.065 165.600 2246.000 166.240 ;
        RECT 4.400 164.200 2246.000 165.600 ;
        RECT 0.065 161.520 2246.000 164.200 ;
        RECT 4.400 160.120 2246.000 161.520 ;
        RECT 0.065 158.120 2246.000 160.120 ;
        RECT 4.400 156.720 2245.600 158.120 ;
        RECT 0.065 154.040 2246.000 156.720 ;
        RECT 4.400 152.640 2246.000 154.040 ;
        RECT 0.065 149.960 2246.000 152.640 ;
        RECT 4.400 148.600 2246.000 149.960 ;
        RECT 4.400 148.560 2245.600 148.600 ;
        RECT 0.065 147.200 2245.600 148.560 ;
        RECT 0.065 146.560 2246.000 147.200 ;
        RECT 4.400 145.160 2246.000 146.560 ;
        RECT 0.065 142.480 2246.000 145.160 ;
        RECT 4.400 141.080 2246.000 142.480 ;
        RECT 0.065 139.080 2246.000 141.080 ;
        RECT 4.400 137.680 2245.600 139.080 ;
        RECT 0.065 135.000 2246.000 137.680 ;
        RECT 4.400 133.600 2246.000 135.000 ;
        RECT 0.065 131.600 2246.000 133.600 ;
        RECT 4.400 130.200 2246.000 131.600 ;
        RECT 0.065 129.560 2246.000 130.200 ;
        RECT 0.065 128.160 2245.600 129.560 ;
        RECT 0.065 127.520 2246.000 128.160 ;
        RECT 4.400 126.120 2246.000 127.520 ;
        RECT 0.065 123.440 2246.000 126.120 ;
        RECT 4.400 122.040 2246.000 123.440 ;
        RECT 0.065 120.040 2246.000 122.040 ;
        RECT 4.400 118.640 2245.600 120.040 ;
        RECT 0.065 115.960 2246.000 118.640 ;
        RECT 4.400 114.560 2246.000 115.960 ;
        RECT 0.065 112.560 2246.000 114.560 ;
        RECT 4.400 111.160 2246.000 112.560 ;
        RECT 0.065 110.520 2246.000 111.160 ;
        RECT 0.065 109.120 2245.600 110.520 ;
        RECT 0.065 108.480 2246.000 109.120 ;
        RECT 4.400 107.080 2246.000 108.480 ;
        RECT 0.065 104.400 2246.000 107.080 ;
        RECT 4.400 103.000 2246.000 104.400 ;
        RECT 0.065 101.000 2246.000 103.000 ;
        RECT 4.400 99.600 2245.600 101.000 ;
        RECT 0.065 96.920 2246.000 99.600 ;
        RECT 4.400 95.520 2246.000 96.920 ;
        RECT 0.065 93.520 2246.000 95.520 ;
        RECT 4.400 92.120 2246.000 93.520 ;
        RECT 0.065 91.480 2246.000 92.120 ;
        RECT 0.065 90.080 2245.600 91.480 ;
        RECT 0.065 89.440 2246.000 90.080 ;
        RECT 4.400 88.040 2246.000 89.440 ;
        RECT 0.065 85.360 2246.000 88.040 ;
        RECT 4.400 83.960 2246.000 85.360 ;
        RECT 0.065 81.960 2246.000 83.960 ;
        RECT 4.400 80.560 2245.600 81.960 ;
        RECT 0.065 77.880 2246.000 80.560 ;
        RECT 4.400 76.480 2246.000 77.880 ;
        RECT 0.065 74.480 2246.000 76.480 ;
        RECT 4.400 73.080 2246.000 74.480 ;
        RECT 0.065 72.440 2246.000 73.080 ;
        RECT 0.065 71.040 2245.600 72.440 ;
        RECT 0.065 70.400 2246.000 71.040 ;
        RECT 4.400 69.000 2246.000 70.400 ;
        RECT 0.065 67.000 2246.000 69.000 ;
        RECT 4.400 65.600 2246.000 67.000 ;
        RECT 0.065 62.920 2246.000 65.600 ;
        RECT 4.400 61.520 2245.600 62.920 ;
        RECT 0.065 58.840 2246.000 61.520 ;
        RECT 4.400 57.440 2246.000 58.840 ;
        RECT 0.065 55.440 2246.000 57.440 ;
        RECT 4.400 54.040 2246.000 55.440 ;
        RECT 0.065 53.400 2246.000 54.040 ;
        RECT 0.065 52.000 2245.600 53.400 ;
        RECT 0.065 51.360 2246.000 52.000 ;
        RECT 4.400 49.960 2246.000 51.360 ;
        RECT 0.065 47.960 2246.000 49.960 ;
        RECT 4.400 46.560 2246.000 47.960 ;
        RECT 0.065 43.880 2246.000 46.560 ;
        RECT 4.400 42.480 2245.600 43.880 ;
        RECT 0.065 39.800 2246.000 42.480 ;
        RECT 4.400 38.400 2246.000 39.800 ;
        RECT 0.065 36.400 2246.000 38.400 ;
        RECT 4.400 35.000 2246.000 36.400 ;
        RECT 0.065 34.360 2246.000 35.000 ;
        RECT 0.065 32.960 2245.600 34.360 ;
        RECT 0.065 32.320 2246.000 32.960 ;
        RECT 4.400 30.920 2246.000 32.320 ;
        RECT 0.065 28.920 2246.000 30.920 ;
        RECT 4.400 27.520 2246.000 28.920 ;
        RECT 0.065 24.840 2246.000 27.520 ;
        RECT 4.400 23.440 2245.600 24.840 ;
        RECT 0.065 20.760 2246.000 23.440 ;
        RECT 4.400 19.360 2246.000 20.760 ;
        RECT 0.065 17.360 2246.000 19.360 ;
        RECT 4.400 15.960 2246.000 17.360 ;
        RECT 0.065 15.320 2246.000 15.960 ;
        RECT 0.065 13.920 2245.600 15.320 ;
        RECT 0.065 13.280 2246.000 13.920 ;
        RECT 4.400 11.880 2246.000 13.280 ;
        RECT 0.065 9.880 2246.000 11.880 ;
        RECT 4.400 8.480 2246.000 9.880 ;
        RECT 0.065 5.800 2246.000 8.480 ;
        RECT 4.400 4.400 2245.600 5.800 ;
        RECT 0.065 2.400 2246.000 4.400 ;
        RECT 4.400 1.540 2246.000 2.400 ;
      LAYER met4 ;
        RECT 9.495 827.520 2234.385 833.505 ;
        RECT 9.495 10.240 20.640 827.520 ;
        RECT 23.040 10.240 45.640 827.520 ;
        RECT 48.040 10.240 70.640 827.520 ;
        RECT 73.040 10.240 95.640 827.520 ;
        RECT 98.040 640.360 120.640 827.520 ;
        RECT 123.040 640.360 145.640 827.520 ;
        RECT 148.040 640.360 170.640 827.520 ;
        RECT 173.040 640.360 195.640 827.520 ;
        RECT 198.040 640.360 220.640 827.520 ;
        RECT 223.040 640.360 245.640 827.520 ;
        RECT 248.040 640.360 270.640 827.520 ;
        RECT 273.040 640.360 295.640 827.520 ;
        RECT 298.040 640.360 320.640 827.520 ;
        RECT 323.040 640.360 345.640 827.520 ;
        RECT 348.040 640.360 370.640 827.520 ;
        RECT 373.040 640.360 395.640 827.520 ;
        RECT 398.040 640.360 420.640 827.520 ;
        RECT 423.040 640.360 445.640 827.520 ;
        RECT 448.040 640.360 470.640 827.520 ;
        RECT 473.040 640.360 495.640 827.520 ;
        RECT 498.040 640.360 520.640 827.520 ;
        RECT 523.040 640.360 545.640 827.520 ;
        RECT 548.040 640.360 570.640 827.520 ;
        RECT 573.040 640.360 595.640 827.520 ;
        RECT 598.040 640.360 620.640 827.520 ;
        RECT 623.040 640.360 645.640 827.520 ;
        RECT 648.040 640.360 670.640 827.520 ;
        RECT 673.040 640.360 695.640 827.520 ;
        RECT 698.040 640.360 720.640 827.520 ;
        RECT 723.040 640.360 745.640 827.520 ;
        RECT 748.040 640.360 770.640 827.520 ;
        RECT 773.040 640.360 795.640 827.520 ;
        RECT 798.040 640.360 820.640 827.520 ;
        RECT 823.040 640.360 845.640 827.520 ;
        RECT 848.040 640.360 870.640 827.520 ;
        RECT 873.040 640.360 895.640 827.520 ;
        RECT 98.040 106.640 895.640 640.360 ;
        RECT 98.040 10.240 120.640 106.640 ;
        RECT 123.040 10.240 145.640 106.640 ;
        RECT 148.040 10.240 170.640 106.640 ;
        RECT 173.040 10.240 195.640 106.640 ;
        RECT 198.040 10.240 220.640 106.640 ;
        RECT 223.040 10.240 245.640 106.640 ;
        RECT 248.040 10.240 270.640 106.640 ;
        RECT 273.040 10.240 295.640 106.640 ;
        RECT 298.040 10.240 320.640 106.640 ;
        RECT 323.040 10.240 345.640 106.640 ;
        RECT 348.040 10.240 370.640 106.640 ;
        RECT 373.040 10.240 395.640 106.640 ;
        RECT 398.040 10.240 420.640 106.640 ;
        RECT 423.040 10.240 445.640 106.640 ;
        RECT 448.040 10.240 470.640 106.640 ;
        RECT 473.040 10.240 495.640 106.640 ;
        RECT 498.040 10.240 520.640 106.640 ;
        RECT 523.040 10.240 545.640 106.640 ;
        RECT 548.040 10.240 570.640 106.640 ;
        RECT 573.040 10.240 595.640 106.640 ;
        RECT 598.040 10.240 620.640 106.640 ;
        RECT 623.040 10.240 645.640 106.640 ;
        RECT 648.040 10.240 670.640 106.640 ;
        RECT 673.040 10.240 695.640 106.640 ;
        RECT 698.040 10.240 720.640 106.640 ;
        RECT 723.040 10.240 745.640 106.640 ;
        RECT 748.040 10.240 770.640 106.640 ;
        RECT 773.040 10.240 795.640 106.640 ;
        RECT 798.040 10.240 820.640 106.640 ;
        RECT 823.040 10.240 845.640 106.640 ;
        RECT 848.040 10.240 870.640 106.640 ;
        RECT 873.040 10.240 895.640 106.640 ;
        RECT 898.040 10.240 920.640 827.520 ;
        RECT 923.040 10.240 945.640 827.520 ;
        RECT 948.040 10.240 970.640 827.520 ;
        RECT 973.040 10.240 995.640 827.520 ;
        RECT 998.040 10.240 1020.640 827.520 ;
        RECT 1023.040 10.240 1045.640 827.520 ;
        RECT 1048.040 10.240 1070.640 827.520 ;
        RECT 1073.040 10.240 1095.640 827.520 ;
        RECT 1098.040 10.240 1120.640 827.520 ;
        RECT 1123.040 10.240 1145.640 827.520 ;
        RECT 1148.040 10.240 1170.640 827.520 ;
        RECT 1173.040 10.240 1195.640 827.520 ;
        RECT 1198.040 10.240 1220.640 827.520 ;
        RECT 1223.040 10.240 1245.640 827.520 ;
        RECT 1248.040 10.240 1270.640 827.520 ;
        RECT 1273.040 10.240 1295.640 827.520 ;
        RECT 1298.040 10.240 1320.640 827.520 ;
        RECT 1323.040 10.240 1345.640 827.520 ;
        RECT 1348.040 10.240 1370.640 827.520 ;
        RECT 1373.040 10.240 1395.640 827.520 ;
        RECT 1398.040 10.240 1420.640 827.520 ;
        RECT 1423.040 10.240 1445.640 827.520 ;
        RECT 1448.040 10.240 1470.640 827.520 ;
        RECT 1473.040 10.240 1495.640 827.520 ;
        RECT 1498.040 10.240 1520.640 827.520 ;
        RECT 1523.040 10.240 1545.640 827.520 ;
        RECT 1548.040 10.240 1570.640 827.520 ;
        RECT 1573.040 10.240 1595.640 827.520 ;
        RECT 1598.040 10.240 1620.640 827.520 ;
        RECT 1623.040 10.240 1645.640 827.520 ;
        RECT 1648.040 10.240 1670.640 827.520 ;
        RECT 1673.040 10.240 1695.640 827.520 ;
        RECT 1698.040 10.240 1720.640 827.520 ;
        RECT 1723.040 10.240 1745.640 827.520 ;
        RECT 1748.040 10.240 1770.640 827.520 ;
        RECT 1773.040 10.240 1795.640 827.520 ;
        RECT 1798.040 10.240 1820.640 827.520 ;
        RECT 1823.040 10.240 1845.640 827.520 ;
        RECT 1848.040 10.240 1870.640 827.520 ;
        RECT 1873.040 10.240 1895.640 827.520 ;
        RECT 1898.040 10.240 1920.640 827.520 ;
        RECT 1923.040 821.080 1945.640 827.520 ;
        RECT 1948.040 821.080 1970.640 827.520 ;
        RECT 1973.040 821.080 1995.640 827.520 ;
        RECT 1998.040 821.080 2020.640 827.520 ;
        RECT 1923.040 727.360 2020.640 821.080 ;
        RECT 1923.040 10.240 1945.640 727.360 ;
        RECT 1948.040 10.240 1970.640 727.360 ;
        RECT 1973.040 10.240 1995.640 727.360 ;
        RECT 1998.040 10.240 2020.640 727.360 ;
        RECT 2023.040 10.240 2045.640 827.520 ;
        RECT 2048.040 10.240 2070.640 827.520 ;
        RECT 2073.040 10.240 2095.640 827.520 ;
        RECT 2098.040 10.240 2120.640 827.520 ;
        RECT 2123.040 10.240 2145.640 827.520 ;
        RECT 2148.040 10.240 2170.640 827.520 ;
        RECT 2173.040 10.240 2195.640 827.520 ;
        RECT 2198.040 10.240 2220.640 827.520 ;
        RECT 2223.040 10.240 2234.385 827.520 ;
        RECT 9.495 1.535 2234.385 10.240 ;
  END
END mgmt_core
END LIBRARY

