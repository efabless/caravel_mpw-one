magic
tech sky130A
magscale 1 2
timestamp 1606509736
<< error_p >>
rect -4395 799 -4337 805
rect -4277 799 -4219 805
rect -4159 799 -4101 805
rect -4041 799 -3983 805
rect -3923 799 -3865 805
rect -3805 799 -3747 805
rect -3687 799 -3629 805
rect -3569 799 -3511 805
rect -3451 799 -3393 805
rect -3333 799 -3275 805
rect -3215 799 -3157 805
rect -3097 799 -3039 805
rect -2979 799 -2921 805
rect -2861 799 -2803 805
rect -2743 799 -2685 805
rect -2625 799 -2567 805
rect -2507 799 -2449 805
rect -2389 799 -2331 805
rect -2271 799 -2213 805
rect -2153 799 -2095 805
rect -2035 799 -1977 805
rect -1917 799 -1859 805
rect -1799 799 -1741 805
rect -1681 799 -1623 805
rect -1563 799 -1505 805
rect -1445 799 -1387 805
rect -1327 799 -1269 805
rect -1209 799 -1151 805
rect -1091 799 -1033 805
rect -973 799 -915 805
rect -855 799 -797 805
rect -737 799 -679 805
rect -619 799 -561 805
rect -501 799 -443 805
rect -383 799 -325 805
rect -265 799 -207 805
rect -147 799 -89 805
rect -29 799 29 805
rect 89 799 147 805
rect 207 799 265 805
rect 325 799 383 805
rect 443 799 501 805
rect 561 799 619 805
rect 679 799 737 805
rect 797 799 855 805
rect 915 799 973 805
rect 1033 799 1091 805
rect 1151 799 1209 805
rect 1269 799 1327 805
rect 1387 799 1445 805
rect 1505 799 1563 805
rect 1623 799 1681 805
rect 1741 799 1799 805
rect 1859 799 1917 805
rect 1977 799 2035 805
rect 2095 799 2153 805
rect 2213 799 2271 805
rect 2331 799 2389 805
rect 2449 799 2507 805
rect 2567 799 2625 805
rect 2685 799 2743 805
rect 2803 799 2861 805
rect 2921 799 2979 805
rect 3039 799 3097 805
rect 3157 799 3215 805
rect 3275 799 3333 805
rect 3393 799 3451 805
rect 3511 799 3569 805
rect 3629 799 3687 805
rect 3747 799 3805 805
rect 3865 799 3923 805
rect 3983 799 4041 805
rect 4101 799 4159 805
rect 4219 799 4277 805
rect 4337 799 4395 805
rect -4395 765 -4383 799
rect -4277 765 -4265 799
rect -4159 765 -4147 799
rect -4041 765 -4029 799
rect -3923 765 -3911 799
rect -3805 765 -3793 799
rect -3687 765 -3675 799
rect -3569 765 -3557 799
rect -3451 765 -3439 799
rect -3333 765 -3321 799
rect -3215 765 -3203 799
rect -3097 765 -3085 799
rect -2979 765 -2967 799
rect -2861 765 -2849 799
rect -2743 765 -2731 799
rect -2625 765 -2613 799
rect -2507 765 -2495 799
rect -2389 765 -2377 799
rect -2271 765 -2259 799
rect -2153 765 -2141 799
rect -2035 765 -2023 799
rect -1917 765 -1905 799
rect -1799 765 -1787 799
rect -1681 765 -1669 799
rect -1563 765 -1551 799
rect -1445 765 -1433 799
rect -1327 765 -1315 799
rect -1209 765 -1197 799
rect -1091 765 -1079 799
rect -973 765 -961 799
rect -855 765 -843 799
rect -737 765 -725 799
rect -619 765 -607 799
rect -501 765 -489 799
rect -383 765 -371 799
rect -265 765 -253 799
rect -147 765 -135 799
rect -29 765 -17 799
rect 89 765 101 799
rect 207 765 219 799
rect 325 765 337 799
rect 443 765 455 799
rect 561 765 573 799
rect 679 765 691 799
rect 797 765 809 799
rect 915 765 927 799
rect 1033 765 1045 799
rect 1151 765 1163 799
rect 1269 765 1281 799
rect 1387 765 1399 799
rect 1505 765 1517 799
rect 1623 765 1635 799
rect 1741 765 1753 799
rect 1859 765 1871 799
rect 1977 765 1989 799
rect 2095 765 2107 799
rect 2213 765 2225 799
rect 2331 765 2343 799
rect 2449 765 2461 799
rect 2567 765 2579 799
rect 2685 765 2697 799
rect 2803 765 2815 799
rect 2921 765 2933 799
rect 3039 765 3051 799
rect 3157 765 3169 799
rect 3275 765 3287 799
rect 3393 765 3405 799
rect 3511 765 3523 799
rect 3629 765 3641 799
rect 3747 765 3759 799
rect 3865 765 3877 799
rect 3983 765 3995 799
rect 4101 765 4113 799
rect 4219 765 4231 799
rect 4337 765 4349 799
rect -4395 759 -4337 765
rect -4277 759 -4219 765
rect -4159 759 -4101 765
rect -4041 759 -3983 765
rect -3923 759 -3865 765
rect -3805 759 -3747 765
rect -3687 759 -3629 765
rect -3569 759 -3511 765
rect -3451 759 -3393 765
rect -3333 759 -3275 765
rect -3215 759 -3157 765
rect -3097 759 -3039 765
rect -2979 759 -2921 765
rect -2861 759 -2803 765
rect -2743 759 -2685 765
rect -2625 759 -2567 765
rect -2507 759 -2449 765
rect -2389 759 -2331 765
rect -2271 759 -2213 765
rect -2153 759 -2095 765
rect -2035 759 -1977 765
rect -1917 759 -1859 765
rect -1799 759 -1741 765
rect -1681 759 -1623 765
rect -1563 759 -1505 765
rect -1445 759 -1387 765
rect -1327 759 -1269 765
rect -1209 759 -1151 765
rect -1091 759 -1033 765
rect -973 759 -915 765
rect -855 759 -797 765
rect -737 759 -679 765
rect -619 759 -561 765
rect -501 759 -443 765
rect -383 759 -325 765
rect -265 759 -207 765
rect -147 759 -89 765
rect -29 759 29 765
rect 89 759 147 765
rect 207 759 265 765
rect 325 759 383 765
rect 443 759 501 765
rect 561 759 619 765
rect 679 759 737 765
rect 797 759 855 765
rect 915 759 973 765
rect 1033 759 1091 765
rect 1151 759 1209 765
rect 1269 759 1327 765
rect 1387 759 1445 765
rect 1505 759 1563 765
rect 1623 759 1681 765
rect 1741 759 1799 765
rect 1859 759 1917 765
rect 1977 759 2035 765
rect 2095 759 2153 765
rect 2213 759 2271 765
rect 2331 759 2389 765
rect 2449 759 2507 765
rect 2567 759 2625 765
rect 2685 759 2743 765
rect 2803 759 2861 765
rect 2921 759 2979 765
rect 3039 759 3097 765
rect 3157 759 3215 765
rect 3275 759 3333 765
rect 3393 759 3451 765
rect 3511 759 3569 765
rect 3629 759 3687 765
rect 3747 759 3805 765
rect 3865 759 3923 765
rect 3983 759 4041 765
rect 4101 759 4159 765
rect 4219 759 4277 765
rect 4337 759 4395 765
rect -4395 71 -4337 77
rect -4277 71 -4219 77
rect -4159 71 -4101 77
rect -4041 71 -3983 77
rect -3923 71 -3865 77
rect -3805 71 -3747 77
rect -3687 71 -3629 77
rect -3569 71 -3511 77
rect -3451 71 -3393 77
rect -3333 71 -3275 77
rect -3215 71 -3157 77
rect -3097 71 -3039 77
rect -2979 71 -2921 77
rect -2861 71 -2803 77
rect -2743 71 -2685 77
rect -2625 71 -2567 77
rect -2507 71 -2449 77
rect -2389 71 -2331 77
rect -2271 71 -2213 77
rect -2153 71 -2095 77
rect -2035 71 -1977 77
rect -1917 71 -1859 77
rect -1799 71 -1741 77
rect -1681 71 -1623 77
rect -1563 71 -1505 77
rect -1445 71 -1387 77
rect -1327 71 -1269 77
rect -1209 71 -1151 77
rect -1091 71 -1033 77
rect -973 71 -915 77
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect 915 71 973 77
rect 1033 71 1091 77
rect 1151 71 1209 77
rect 1269 71 1327 77
rect 1387 71 1445 77
rect 1505 71 1563 77
rect 1623 71 1681 77
rect 1741 71 1799 77
rect 1859 71 1917 77
rect 1977 71 2035 77
rect 2095 71 2153 77
rect 2213 71 2271 77
rect 2331 71 2389 77
rect 2449 71 2507 77
rect 2567 71 2625 77
rect 2685 71 2743 77
rect 2803 71 2861 77
rect 2921 71 2979 77
rect 3039 71 3097 77
rect 3157 71 3215 77
rect 3275 71 3333 77
rect 3393 71 3451 77
rect 3511 71 3569 77
rect 3629 71 3687 77
rect 3747 71 3805 77
rect 3865 71 3923 77
rect 3983 71 4041 77
rect 4101 71 4159 77
rect 4219 71 4277 77
rect 4337 71 4395 77
rect -4395 37 -4383 71
rect -4277 37 -4265 71
rect -4159 37 -4147 71
rect -4041 37 -4029 71
rect -3923 37 -3911 71
rect -3805 37 -3793 71
rect -3687 37 -3675 71
rect -3569 37 -3557 71
rect -3451 37 -3439 71
rect -3333 37 -3321 71
rect -3215 37 -3203 71
rect -3097 37 -3085 71
rect -2979 37 -2967 71
rect -2861 37 -2849 71
rect -2743 37 -2731 71
rect -2625 37 -2613 71
rect -2507 37 -2495 71
rect -2389 37 -2377 71
rect -2271 37 -2259 71
rect -2153 37 -2141 71
rect -2035 37 -2023 71
rect -1917 37 -1905 71
rect -1799 37 -1787 71
rect -1681 37 -1669 71
rect -1563 37 -1551 71
rect -1445 37 -1433 71
rect -1327 37 -1315 71
rect -1209 37 -1197 71
rect -1091 37 -1079 71
rect -973 37 -961 71
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect 915 37 927 71
rect 1033 37 1045 71
rect 1151 37 1163 71
rect 1269 37 1281 71
rect 1387 37 1399 71
rect 1505 37 1517 71
rect 1623 37 1635 71
rect 1741 37 1753 71
rect 1859 37 1871 71
rect 1977 37 1989 71
rect 2095 37 2107 71
rect 2213 37 2225 71
rect 2331 37 2343 71
rect 2449 37 2461 71
rect 2567 37 2579 71
rect 2685 37 2697 71
rect 2803 37 2815 71
rect 2921 37 2933 71
rect 3039 37 3051 71
rect 3157 37 3169 71
rect 3275 37 3287 71
rect 3393 37 3405 71
rect 3511 37 3523 71
rect 3629 37 3641 71
rect 3747 37 3759 71
rect 3865 37 3877 71
rect 3983 37 3995 71
rect 4101 37 4113 71
rect 4219 37 4231 71
rect 4337 37 4349 71
rect -4395 31 -4337 37
rect -4277 31 -4219 37
rect -4159 31 -4101 37
rect -4041 31 -3983 37
rect -3923 31 -3865 37
rect -3805 31 -3747 37
rect -3687 31 -3629 37
rect -3569 31 -3511 37
rect -3451 31 -3393 37
rect -3333 31 -3275 37
rect -3215 31 -3157 37
rect -3097 31 -3039 37
rect -2979 31 -2921 37
rect -2861 31 -2803 37
rect -2743 31 -2685 37
rect -2625 31 -2567 37
rect -2507 31 -2449 37
rect -2389 31 -2331 37
rect -2271 31 -2213 37
rect -2153 31 -2095 37
rect -2035 31 -1977 37
rect -1917 31 -1859 37
rect -1799 31 -1741 37
rect -1681 31 -1623 37
rect -1563 31 -1505 37
rect -1445 31 -1387 37
rect -1327 31 -1269 37
rect -1209 31 -1151 37
rect -1091 31 -1033 37
rect -973 31 -915 37
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect 915 31 973 37
rect 1033 31 1091 37
rect 1151 31 1209 37
rect 1269 31 1327 37
rect 1387 31 1445 37
rect 1505 31 1563 37
rect 1623 31 1681 37
rect 1741 31 1799 37
rect 1859 31 1917 37
rect 1977 31 2035 37
rect 2095 31 2153 37
rect 2213 31 2271 37
rect 2331 31 2389 37
rect 2449 31 2507 37
rect 2567 31 2625 37
rect 2685 31 2743 37
rect 2803 31 2861 37
rect 2921 31 2979 37
rect 3039 31 3097 37
rect 3157 31 3215 37
rect 3275 31 3333 37
rect 3393 31 3451 37
rect 3511 31 3569 37
rect 3629 31 3687 37
rect 3747 31 3805 37
rect 3865 31 3923 37
rect 3983 31 4041 37
rect 4101 31 4159 37
rect 4219 31 4277 37
rect 4337 31 4395 37
rect -4395 -37 -4337 -31
rect -4277 -37 -4219 -31
rect -4159 -37 -4101 -31
rect -4041 -37 -3983 -31
rect -3923 -37 -3865 -31
rect -3805 -37 -3747 -31
rect -3687 -37 -3629 -31
rect -3569 -37 -3511 -31
rect -3451 -37 -3393 -31
rect -3333 -37 -3275 -31
rect -3215 -37 -3157 -31
rect -3097 -37 -3039 -31
rect -2979 -37 -2921 -31
rect -2861 -37 -2803 -31
rect -2743 -37 -2685 -31
rect -2625 -37 -2567 -31
rect -2507 -37 -2449 -31
rect -2389 -37 -2331 -31
rect -2271 -37 -2213 -31
rect -2153 -37 -2095 -31
rect -2035 -37 -1977 -31
rect -1917 -37 -1859 -31
rect -1799 -37 -1741 -31
rect -1681 -37 -1623 -31
rect -1563 -37 -1505 -31
rect -1445 -37 -1387 -31
rect -1327 -37 -1269 -31
rect -1209 -37 -1151 -31
rect -1091 -37 -1033 -31
rect -973 -37 -915 -31
rect -855 -37 -797 -31
rect -737 -37 -679 -31
rect -619 -37 -561 -31
rect -501 -37 -443 -31
rect -383 -37 -325 -31
rect -265 -37 -207 -31
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect 207 -37 265 -31
rect 325 -37 383 -31
rect 443 -37 501 -31
rect 561 -37 619 -31
rect 679 -37 737 -31
rect 797 -37 855 -31
rect 915 -37 973 -31
rect 1033 -37 1091 -31
rect 1151 -37 1209 -31
rect 1269 -37 1327 -31
rect 1387 -37 1445 -31
rect 1505 -37 1563 -31
rect 1623 -37 1681 -31
rect 1741 -37 1799 -31
rect 1859 -37 1917 -31
rect 1977 -37 2035 -31
rect 2095 -37 2153 -31
rect 2213 -37 2271 -31
rect 2331 -37 2389 -31
rect 2449 -37 2507 -31
rect 2567 -37 2625 -31
rect 2685 -37 2743 -31
rect 2803 -37 2861 -31
rect 2921 -37 2979 -31
rect 3039 -37 3097 -31
rect 3157 -37 3215 -31
rect 3275 -37 3333 -31
rect 3393 -37 3451 -31
rect 3511 -37 3569 -31
rect 3629 -37 3687 -31
rect 3747 -37 3805 -31
rect 3865 -37 3923 -31
rect 3983 -37 4041 -31
rect 4101 -37 4159 -31
rect 4219 -37 4277 -31
rect 4337 -37 4395 -31
rect -4395 -71 -4383 -37
rect -4277 -71 -4265 -37
rect -4159 -71 -4147 -37
rect -4041 -71 -4029 -37
rect -3923 -71 -3911 -37
rect -3805 -71 -3793 -37
rect -3687 -71 -3675 -37
rect -3569 -71 -3557 -37
rect -3451 -71 -3439 -37
rect -3333 -71 -3321 -37
rect -3215 -71 -3203 -37
rect -3097 -71 -3085 -37
rect -2979 -71 -2967 -37
rect -2861 -71 -2849 -37
rect -2743 -71 -2731 -37
rect -2625 -71 -2613 -37
rect -2507 -71 -2495 -37
rect -2389 -71 -2377 -37
rect -2271 -71 -2259 -37
rect -2153 -71 -2141 -37
rect -2035 -71 -2023 -37
rect -1917 -71 -1905 -37
rect -1799 -71 -1787 -37
rect -1681 -71 -1669 -37
rect -1563 -71 -1551 -37
rect -1445 -71 -1433 -37
rect -1327 -71 -1315 -37
rect -1209 -71 -1197 -37
rect -1091 -71 -1079 -37
rect -973 -71 -961 -37
rect -855 -71 -843 -37
rect -737 -71 -725 -37
rect -619 -71 -607 -37
rect -501 -71 -489 -37
rect -383 -71 -371 -37
rect -265 -71 -253 -37
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect 207 -71 219 -37
rect 325 -71 337 -37
rect 443 -71 455 -37
rect 561 -71 573 -37
rect 679 -71 691 -37
rect 797 -71 809 -37
rect 915 -71 927 -37
rect 1033 -71 1045 -37
rect 1151 -71 1163 -37
rect 1269 -71 1281 -37
rect 1387 -71 1399 -37
rect 1505 -71 1517 -37
rect 1623 -71 1635 -37
rect 1741 -71 1753 -37
rect 1859 -71 1871 -37
rect 1977 -71 1989 -37
rect 2095 -71 2107 -37
rect 2213 -71 2225 -37
rect 2331 -71 2343 -37
rect 2449 -71 2461 -37
rect 2567 -71 2579 -37
rect 2685 -71 2697 -37
rect 2803 -71 2815 -37
rect 2921 -71 2933 -37
rect 3039 -71 3051 -37
rect 3157 -71 3169 -37
rect 3275 -71 3287 -37
rect 3393 -71 3405 -37
rect 3511 -71 3523 -37
rect 3629 -71 3641 -37
rect 3747 -71 3759 -37
rect 3865 -71 3877 -37
rect 3983 -71 3995 -37
rect 4101 -71 4113 -37
rect 4219 -71 4231 -37
rect 4337 -71 4349 -37
rect -4395 -77 -4337 -71
rect -4277 -77 -4219 -71
rect -4159 -77 -4101 -71
rect -4041 -77 -3983 -71
rect -3923 -77 -3865 -71
rect -3805 -77 -3747 -71
rect -3687 -77 -3629 -71
rect -3569 -77 -3511 -71
rect -3451 -77 -3393 -71
rect -3333 -77 -3275 -71
rect -3215 -77 -3157 -71
rect -3097 -77 -3039 -71
rect -2979 -77 -2921 -71
rect -2861 -77 -2803 -71
rect -2743 -77 -2685 -71
rect -2625 -77 -2567 -71
rect -2507 -77 -2449 -71
rect -2389 -77 -2331 -71
rect -2271 -77 -2213 -71
rect -2153 -77 -2095 -71
rect -2035 -77 -1977 -71
rect -1917 -77 -1859 -71
rect -1799 -77 -1741 -71
rect -1681 -77 -1623 -71
rect -1563 -77 -1505 -71
rect -1445 -77 -1387 -71
rect -1327 -77 -1269 -71
rect -1209 -77 -1151 -71
rect -1091 -77 -1033 -71
rect -973 -77 -915 -71
rect -855 -77 -797 -71
rect -737 -77 -679 -71
rect -619 -77 -561 -71
rect -501 -77 -443 -71
rect -383 -77 -325 -71
rect -265 -77 -207 -71
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect 207 -77 265 -71
rect 325 -77 383 -71
rect 443 -77 501 -71
rect 561 -77 619 -71
rect 679 -77 737 -71
rect 797 -77 855 -71
rect 915 -77 973 -71
rect 1033 -77 1091 -71
rect 1151 -77 1209 -71
rect 1269 -77 1327 -71
rect 1387 -77 1445 -71
rect 1505 -77 1563 -71
rect 1623 -77 1681 -71
rect 1741 -77 1799 -71
rect 1859 -77 1917 -71
rect 1977 -77 2035 -71
rect 2095 -77 2153 -71
rect 2213 -77 2271 -71
rect 2331 -77 2389 -71
rect 2449 -77 2507 -71
rect 2567 -77 2625 -71
rect 2685 -77 2743 -71
rect 2803 -77 2861 -71
rect 2921 -77 2979 -71
rect 3039 -77 3097 -71
rect 3157 -77 3215 -71
rect 3275 -77 3333 -71
rect 3393 -77 3451 -71
rect 3511 -77 3569 -71
rect 3629 -77 3687 -71
rect 3747 -77 3805 -71
rect 3865 -77 3923 -71
rect 3983 -77 4041 -71
rect 4101 -77 4159 -71
rect 4219 -77 4277 -71
rect 4337 -77 4395 -71
rect -4395 -765 -4337 -759
rect -4277 -765 -4219 -759
rect -4159 -765 -4101 -759
rect -4041 -765 -3983 -759
rect -3923 -765 -3865 -759
rect -3805 -765 -3747 -759
rect -3687 -765 -3629 -759
rect -3569 -765 -3511 -759
rect -3451 -765 -3393 -759
rect -3333 -765 -3275 -759
rect -3215 -765 -3157 -759
rect -3097 -765 -3039 -759
rect -2979 -765 -2921 -759
rect -2861 -765 -2803 -759
rect -2743 -765 -2685 -759
rect -2625 -765 -2567 -759
rect -2507 -765 -2449 -759
rect -2389 -765 -2331 -759
rect -2271 -765 -2213 -759
rect -2153 -765 -2095 -759
rect -2035 -765 -1977 -759
rect -1917 -765 -1859 -759
rect -1799 -765 -1741 -759
rect -1681 -765 -1623 -759
rect -1563 -765 -1505 -759
rect -1445 -765 -1387 -759
rect -1327 -765 -1269 -759
rect -1209 -765 -1151 -759
rect -1091 -765 -1033 -759
rect -973 -765 -915 -759
rect -855 -765 -797 -759
rect -737 -765 -679 -759
rect -619 -765 -561 -759
rect -501 -765 -443 -759
rect -383 -765 -325 -759
rect -265 -765 -207 -759
rect -147 -765 -89 -759
rect -29 -765 29 -759
rect 89 -765 147 -759
rect 207 -765 265 -759
rect 325 -765 383 -759
rect 443 -765 501 -759
rect 561 -765 619 -759
rect 679 -765 737 -759
rect 797 -765 855 -759
rect 915 -765 973 -759
rect 1033 -765 1091 -759
rect 1151 -765 1209 -759
rect 1269 -765 1327 -759
rect 1387 -765 1445 -759
rect 1505 -765 1563 -759
rect 1623 -765 1681 -759
rect 1741 -765 1799 -759
rect 1859 -765 1917 -759
rect 1977 -765 2035 -759
rect 2095 -765 2153 -759
rect 2213 -765 2271 -759
rect 2331 -765 2389 -759
rect 2449 -765 2507 -759
rect 2567 -765 2625 -759
rect 2685 -765 2743 -759
rect 2803 -765 2861 -759
rect 2921 -765 2979 -759
rect 3039 -765 3097 -759
rect 3157 -765 3215 -759
rect 3275 -765 3333 -759
rect 3393 -765 3451 -759
rect 3511 -765 3569 -759
rect 3629 -765 3687 -759
rect 3747 -765 3805 -759
rect 3865 -765 3923 -759
rect 3983 -765 4041 -759
rect 4101 -765 4159 -759
rect 4219 -765 4277 -759
rect 4337 -765 4395 -759
rect -4395 -799 -4383 -765
rect -4277 -799 -4265 -765
rect -4159 -799 -4147 -765
rect -4041 -799 -4029 -765
rect -3923 -799 -3911 -765
rect -3805 -799 -3793 -765
rect -3687 -799 -3675 -765
rect -3569 -799 -3557 -765
rect -3451 -799 -3439 -765
rect -3333 -799 -3321 -765
rect -3215 -799 -3203 -765
rect -3097 -799 -3085 -765
rect -2979 -799 -2967 -765
rect -2861 -799 -2849 -765
rect -2743 -799 -2731 -765
rect -2625 -799 -2613 -765
rect -2507 -799 -2495 -765
rect -2389 -799 -2377 -765
rect -2271 -799 -2259 -765
rect -2153 -799 -2141 -765
rect -2035 -799 -2023 -765
rect -1917 -799 -1905 -765
rect -1799 -799 -1787 -765
rect -1681 -799 -1669 -765
rect -1563 -799 -1551 -765
rect -1445 -799 -1433 -765
rect -1327 -799 -1315 -765
rect -1209 -799 -1197 -765
rect -1091 -799 -1079 -765
rect -973 -799 -961 -765
rect -855 -799 -843 -765
rect -737 -799 -725 -765
rect -619 -799 -607 -765
rect -501 -799 -489 -765
rect -383 -799 -371 -765
rect -265 -799 -253 -765
rect -147 -799 -135 -765
rect -29 -799 -17 -765
rect 89 -799 101 -765
rect 207 -799 219 -765
rect 325 -799 337 -765
rect 443 -799 455 -765
rect 561 -799 573 -765
rect 679 -799 691 -765
rect 797 -799 809 -765
rect 915 -799 927 -765
rect 1033 -799 1045 -765
rect 1151 -799 1163 -765
rect 1269 -799 1281 -765
rect 1387 -799 1399 -765
rect 1505 -799 1517 -765
rect 1623 -799 1635 -765
rect 1741 -799 1753 -765
rect 1859 -799 1871 -765
rect 1977 -799 1989 -765
rect 2095 -799 2107 -765
rect 2213 -799 2225 -765
rect 2331 -799 2343 -765
rect 2449 -799 2461 -765
rect 2567 -799 2579 -765
rect 2685 -799 2697 -765
rect 2803 -799 2815 -765
rect 2921 -799 2933 -765
rect 3039 -799 3051 -765
rect 3157 -799 3169 -765
rect 3275 -799 3287 -765
rect 3393 -799 3405 -765
rect 3511 -799 3523 -765
rect 3629 -799 3641 -765
rect 3747 -799 3759 -765
rect 3865 -799 3877 -765
rect 3983 -799 3995 -765
rect 4101 -799 4113 -765
rect 4219 -799 4231 -765
rect 4337 -799 4349 -765
rect -4395 -805 -4337 -799
rect -4277 -805 -4219 -799
rect -4159 -805 -4101 -799
rect -4041 -805 -3983 -799
rect -3923 -805 -3865 -799
rect -3805 -805 -3747 -799
rect -3687 -805 -3629 -799
rect -3569 -805 -3511 -799
rect -3451 -805 -3393 -799
rect -3333 -805 -3275 -799
rect -3215 -805 -3157 -799
rect -3097 -805 -3039 -799
rect -2979 -805 -2921 -799
rect -2861 -805 -2803 -799
rect -2743 -805 -2685 -799
rect -2625 -805 -2567 -799
rect -2507 -805 -2449 -799
rect -2389 -805 -2331 -799
rect -2271 -805 -2213 -799
rect -2153 -805 -2095 -799
rect -2035 -805 -1977 -799
rect -1917 -805 -1859 -799
rect -1799 -805 -1741 -799
rect -1681 -805 -1623 -799
rect -1563 -805 -1505 -799
rect -1445 -805 -1387 -799
rect -1327 -805 -1269 -799
rect -1209 -805 -1151 -799
rect -1091 -805 -1033 -799
rect -973 -805 -915 -799
rect -855 -805 -797 -799
rect -737 -805 -679 -799
rect -619 -805 -561 -799
rect -501 -805 -443 -799
rect -383 -805 -325 -799
rect -265 -805 -207 -799
rect -147 -805 -89 -799
rect -29 -805 29 -799
rect 89 -805 147 -799
rect 207 -805 265 -799
rect 325 -805 383 -799
rect 443 -805 501 -799
rect 561 -805 619 -799
rect 679 -805 737 -799
rect 797 -805 855 -799
rect 915 -805 973 -799
rect 1033 -805 1091 -799
rect 1151 -805 1209 -799
rect 1269 -805 1327 -799
rect 1387 -805 1445 -799
rect 1505 -805 1563 -799
rect 1623 -805 1681 -799
rect 1741 -805 1799 -799
rect 1859 -805 1917 -799
rect 1977 -805 2035 -799
rect 2095 -805 2153 -799
rect 2213 -805 2271 -799
rect 2331 -805 2389 -799
rect 2449 -805 2507 -799
rect 2567 -805 2625 -799
rect 2685 -805 2743 -799
rect 2803 -805 2861 -799
rect 2921 -805 2979 -799
rect 3039 -805 3097 -799
rect 3157 -805 3215 -799
rect 3275 -805 3333 -799
rect 3393 -805 3451 -799
rect 3511 -805 3569 -799
rect 3629 -805 3687 -799
rect 3747 -805 3805 -799
rect 3865 -805 3923 -799
rect 3983 -805 4041 -799
rect 4101 -805 4159 -799
rect 4219 -805 4277 -799
rect 4337 -805 4395 -799
<< nwell >>
rect -4592 -937 4592 937
<< pmos >>
rect -4396 118 -4336 718
rect -4278 118 -4218 718
rect -4160 118 -4100 718
rect -4042 118 -3982 718
rect -3924 118 -3864 718
rect -3806 118 -3746 718
rect -3688 118 -3628 718
rect -3570 118 -3510 718
rect -3452 118 -3392 718
rect -3334 118 -3274 718
rect -3216 118 -3156 718
rect -3098 118 -3038 718
rect -2980 118 -2920 718
rect -2862 118 -2802 718
rect -2744 118 -2684 718
rect -2626 118 -2566 718
rect -2508 118 -2448 718
rect -2390 118 -2330 718
rect -2272 118 -2212 718
rect -2154 118 -2094 718
rect -2036 118 -1976 718
rect -1918 118 -1858 718
rect -1800 118 -1740 718
rect -1682 118 -1622 718
rect -1564 118 -1504 718
rect -1446 118 -1386 718
rect -1328 118 -1268 718
rect -1210 118 -1150 718
rect -1092 118 -1032 718
rect -974 118 -914 718
rect -856 118 -796 718
rect -738 118 -678 718
rect -620 118 -560 718
rect -502 118 -442 718
rect -384 118 -324 718
rect -266 118 -206 718
rect -148 118 -88 718
rect -30 118 30 718
rect 88 118 148 718
rect 206 118 266 718
rect 324 118 384 718
rect 442 118 502 718
rect 560 118 620 718
rect 678 118 738 718
rect 796 118 856 718
rect 914 118 974 718
rect 1032 118 1092 718
rect 1150 118 1210 718
rect 1268 118 1328 718
rect 1386 118 1446 718
rect 1504 118 1564 718
rect 1622 118 1682 718
rect 1740 118 1800 718
rect 1858 118 1918 718
rect 1976 118 2036 718
rect 2094 118 2154 718
rect 2212 118 2272 718
rect 2330 118 2390 718
rect 2448 118 2508 718
rect 2566 118 2626 718
rect 2684 118 2744 718
rect 2802 118 2862 718
rect 2920 118 2980 718
rect 3038 118 3098 718
rect 3156 118 3216 718
rect 3274 118 3334 718
rect 3392 118 3452 718
rect 3510 118 3570 718
rect 3628 118 3688 718
rect 3746 118 3806 718
rect 3864 118 3924 718
rect 3982 118 4042 718
rect 4100 118 4160 718
rect 4218 118 4278 718
rect 4336 118 4396 718
rect -4396 -718 -4336 -118
rect -4278 -718 -4218 -118
rect -4160 -718 -4100 -118
rect -4042 -718 -3982 -118
rect -3924 -718 -3864 -118
rect -3806 -718 -3746 -118
rect -3688 -718 -3628 -118
rect -3570 -718 -3510 -118
rect -3452 -718 -3392 -118
rect -3334 -718 -3274 -118
rect -3216 -718 -3156 -118
rect -3098 -718 -3038 -118
rect -2980 -718 -2920 -118
rect -2862 -718 -2802 -118
rect -2744 -718 -2684 -118
rect -2626 -718 -2566 -118
rect -2508 -718 -2448 -118
rect -2390 -718 -2330 -118
rect -2272 -718 -2212 -118
rect -2154 -718 -2094 -118
rect -2036 -718 -1976 -118
rect -1918 -718 -1858 -118
rect -1800 -718 -1740 -118
rect -1682 -718 -1622 -118
rect -1564 -718 -1504 -118
rect -1446 -718 -1386 -118
rect -1328 -718 -1268 -118
rect -1210 -718 -1150 -118
rect -1092 -718 -1032 -118
rect -974 -718 -914 -118
rect -856 -718 -796 -118
rect -738 -718 -678 -118
rect -620 -718 -560 -118
rect -502 -718 -442 -118
rect -384 -718 -324 -118
rect -266 -718 -206 -118
rect -148 -718 -88 -118
rect -30 -718 30 -118
rect 88 -718 148 -118
rect 206 -718 266 -118
rect 324 -718 384 -118
rect 442 -718 502 -118
rect 560 -718 620 -118
rect 678 -718 738 -118
rect 796 -718 856 -118
rect 914 -718 974 -118
rect 1032 -718 1092 -118
rect 1150 -718 1210 -118
rect 1268 -718 1328 -118
rect 1386 -718 1446 -118
rect 1504 -718 1564 -118
rect 1622 -718 1682 -118
rect 1740 -718 1800 -118
rect 1858 -718 1918 -118
rect 1976 -718 2036 -118
rect 2094 -718 2154 -118
rect 2212 -718 2272 -118
rect 2330 -718 2390 -118
rect 2448 -718 2508 -118
rect 2566 -718 2626 -118
rect 2684 -718 2744 -118
rect 2802 -718 2862 -118
rect 2920 -718 2980 -118
rect 3038 -718 3098 -118
rect 3156 -718 3216 -118
rect 3274 -718 3334 -118
rect 3392 -718 3452 -118
rect 3510 -718 3570 -118
rect 3628 -718 3688 -118
rect 3746 -718 3806 -118
rect 3864 -718 3924 -118
rect 3982 -718 4042 -118
rect 4100 -718 4160 -118
rect 4218 -718 4278 -118
rect 4336 -718 4396 -118
<< pdiff >>
rect -4454 706 -4396 718
rect -4454 130 -4442 706
rect -4408 130 -4396 706
rect -4454 118 -4396 130
rect -4336 706 -4278 718
rect -4336 130 -4324 706
rect -4290 130 -4278 706
rect -4336 118 -4278 130
rect -4218 706 -4160 718
rect -4218 130 -4206 706
rect -4172 130 -4160 706
rect -4218 118 -4160 130
rect -4100 706 -4042 718
rect -4100 130 -4088 706
rect -4054 130 -4042 706
rect -4100 118 -4042 130
rect -3982 706 -3924 718
rect -3982 130 -3970 706
rect -3936 130 -3924 706
rect -3982 118 -3924 130
rect -3864 706 -3806 718
rect -3864 130 -3852 706
rect -3818 130 -3806 706
rect -3864 118 -3806 130
rect -3746 706 -3688 718
rect -3746 130 -3734 706
rect -3700 130 -3688 706
rect -3746 118 -3688 130
rect -3628 706 -3570 718
rect -3628 130 -3616 706
rect -3582 130 -3570 706
rect -3628 118 -3570 130
rect -3510 706 -3452 718
rect -3510 130 -3498 706
rect -3464 130 -3452 706
rect -3510 118 -3452 130
rect -3392 706 -3334 718
rect -3392 130 -3380 706
rect -3346 130 -3334 706
rect -3392 118 -3334 130
rect -3274 706 -3216 718
rect -3274 130 -3262 706
rect -3228 130 -3216 706
rect -3274 118 -3216 130
rect -3156 706 -3098 718
rect -3156 130 -3144 706
rect -3110 130 -3098 706
rect -3156 118 -3098 130
rect -3038 706 -2980 718
rect -3038 130 -3026 706
rect -2992 130 -2980 706
rect -3038 118 -2980 130
rect -2920 706 -2862 718
rect -2920 130 -2908 706
rect -2874 130 -2862 706
rect -2920 118 -2862 130
rect -2802 706 -2744 718
rect -2802 130 -2790 706
rect -2756 130 -2744 706
rect -2802 118 -2744 130
rect -2684 706 -2626 718
rect -2684 130 -2672 706
rect -2638 130 -2626 706
rect -2684 118 -2626 130
rect -2566 706 -2508 718
rect -2566 130 -2554 706
rect -2520 130 -2508 706
rect -2566 118 -2508 130
rect -2448 706 -2390 718
rect -2448 130 -2436 706
rect -2402 130 -2390 706
rect -2448 118 -2390 130
rect -2330 706 -2272 718
rect -2330 130 -2318 706
rect -2284 130 -2272 706
rect -2330 118 -2272 130
rect -2212 706 -2154 718
rect -2212 130 -2200 706
rect -2166 130 -2154 706
rect -2212 118 -2154 130
rect -2094 706 -2036 718
rect -2094 130 -2082 706
rect -2048 130 -2036 706
rect -2094 118 -2036 130
rect -1976 706 -1918 718
rect -1976 130 -1964 706
rect -1930 130 -1918 706
rect -1976 118 -1918 130
rect -1858 706 -1800 718
rect -1858 130 -1846 706
rect -1812 130 -1800 706
rect -1858 118 -1800 130
rect -1740 706 -1682 718
rect -1740 130 -1728 706
rect -1694 130 -1682 706
rect -1740 118 -1682 130
rect -1622 706 -1564 718
rect -1622 130 -1610 706
rect -1576 130 -1564 706
rect -1622 118 -1564 130
rect -1504 706 -1446 718
rect -1504 130 -1492 706
rect -1458 130 -1446 706
rect -1504 118 -1446 130
rect -1386 706 -1328 718
rect -1386 130 -1374 706
rect -1340 130 -1328 706
rect -1386 118 -1328 130
rect -1268 706 -1210 718
rect -1268 130 -1256 706
rect -1222 130 -1210 706
rect -1268 118 -1210 130
rect -1150 706 -1092 718
rect -1150 130 -1138 706
rect -1104 130 -1092 706
rect -1150 118 -1092 130
rect -1032 706 -974 718
rect -1032 130 -1020 706
rect -986 130 -974 706
rect -1032 118 -974 130
rect -914 706 -856 718
rect -914 130 -902 706
rect -868 130 -856 706
rect -914 118 -856 130
rect -796 706 -738 718
rect -796 130 -784 706
rect -750 130 -738 706
rect -796 118 -738 130
rect -678 706 -620 718
rect -678 130 -666 706
rect -632 130 -620 706
rect -678 118 -620 130
rect -560 706 -502 718
rect -560 130 -548 706
rect -514 130 -502 706
rect -560 118 -502 130
rect -442 706 -384 718
rect -442 130 -430 706
rect -396 130 -384 706
rect -442 118 -384 130
rect -324 706 -266 718
rect -324 130 -312 706
rect -278 130 -266 706
rect -324 118 -266 130
rect -206 706 -148 718
rect -206 130 -194 706
rect -160 130 -148 706
rect -206 118 -148 130
rect -88 706 -30 718
rect -88 130 -76 706
rect -42 130 -30 706
rect -88 118 -30 130
rect 30 706 88 718
rect 30 130 42 706
rect 76 130 88 706
rect 30 118 88 130
rect 148 706 206 718
rect 148 130 160 706
rect 194 130 206 706
rect 148 118 206 130
rect 266 706 324 718
rect 266 130 278 706
rect 312 130 324 706
rect 266 118 324 130
rect 384 706 442 718
rect 384 130 396 706
rect 430 130 442 706
rect 384 118 442 130
rect 502 706 560 718
rect 502 130 514 706
rect 548 130 560 706
rect 502 118 560 130
rect 620 706 678 718
rect 620 130 632 706
rect 666 130 678 706
rect 620 118 678 130
rect 738 706 796 718
rect 738 130 750 706
rect 784 130 796 706
rect 738 118 796 130
rect 856 706 914 718
rect 856 130 868 706
rect 902 130 914 706
rect 856 118 914 130
rect 974 706 1032 718
rect 974 130 986 706
rect 1020 130 1032 706
rect 974 118 1032 130
rect 1092 706 1150 718
rect 1092 130 1104 706
rect 1138 130 1150 706
rect 1092 118 1150 130
rect 1210 706 1268 718
rect 1210 130 1222 706
rect 1256 130 1268 706
rect 1210 118 1268 130
rect 1328 706 1386 718
rect 1328 130 1340 706
rect 1374 130 1386 706
rect 1328 118 1386 130
rect 1446 706 1504 718
rect 1446 130 1458 706
rect 1492 130 1504 706
rect 1446 118 1504 130
rect 1564 706 1622 718
rect 1564 130 1576 706
rect 1610 130 1622 706
rect 1564 118 1622 130
rect 1682 706 1740 718
rect 1682 130 1694 706
rect 1728 130 1740 706
rect 1682 118 1740 130
rect 1800 706 1858 718
rect 1800 130 1812 706
rect 1846 130 1858 706
rect 1800 118 1858 130
rect 1918 706 1976 718
rect 1918 130 1930 706
rect 1964 130 1976 706
rect 1918 118 1976 130
rect 2036 706 2094 718
rect 2036 130 2048 706
rect 2082 130 2094 706
rect 2036 118 2094 130
rect 2154 706 2212 718
rect 2154 130 2166 706
rect 2200 130 2212 706
rect 2154 118 2212 130
rect 2272 706 2330 718
rect 2272 130 2284 706
rect 2318 130 2330 706
rect 2272 118 2330 130
rect 2390 706 2448 718
rect 2390 130 2402 706
rect 2436 130 2448 706
rect 2390 118 2448 130
rect 2508 706 2566 718
rect 2508 130 2520 706
rect 2554 130 2566 706
rect 2508 118 2566 130
rect 2626 706 2684 718
rect 2626 130 2638 706
rect 2672 130 2684 706
rect 2626 118 2684 130
rect 2744 706 2802 718
rect 2744 130 2756 706
rect 2790 130 2802 706
rect 2744 118 2802 130
rect 2862 706 2920 718
rect 2862 130 2874 706
rect 2908 130 2920 706
rect 2862 118 2920 130
rect 2980 706 3038 718
rect 2980 130 2992 706
rect 3026 130 3038 706
rect 2980 118 3038 130
rect 3098 706 3156 718
rect 3098 130 3110 706
rect 3144 130 3156 706
rect 3098 118 3156 130
rect 3216 706 3274 718
rect 3216 130 3228 706
rect 3262 130 3274 706
rect 3216 118 3274 130
rect 3334 706 3392 718
rect 3334 130 3346 706
rect 3380 130 3392 706
rect 3334 118 3392 130
rect 3452 706 3510 718
rect 3452 130 3464 706
rect 3498 130 3510 706
rect 3452 118 3510 130
rect 3570 706 3628 718
rect 3570 130 3582 706
rect 3616 130 3628 706
rect 3570 118 3628 130
rect 3688 706 3746 718
rect 3688 130 3700 706
rect 3734 130 3746 706
rect 3688 118 3746 130
rect 3806 706 3864 718
rect 3806 130 3818 706
rect 3852 130 3864 706
rect 3806 118 3864 130
rect 3924 706 3982 718
rect 3924 130 3936 706
rect 3970 130 3982 706
rect 3924 118 3982 130
rect 4042 706 4100 718
rect 4042 130 4054 706
rect 4088 130 4100 706
rect 4042 118 4100 130
rect 4160 706 4218 718
rect 4160 130 4172 706
rect 4206 130 4218 706
rect 4160 118 4218 130
rect 4278 706 4336 718
rect 4278 130 4290 706
rect 4324 130 4336 706
rect 4278 118 4336 130
rect 4396 706 4454 718
rect 4396 130 4408 706
rect 4442 130 4454 706
rect 4396 118 4454 130
rect -4454 -130 -4396 -118
rect -4454 -706 -4442 -130
rect -4408 -706 -4396 -130
rect -4454 -718 -4396 -706
rect -4336 -130 -4278 -118
rect -4336 -706 -4324 -130
rect -4290 -706 -4278 -130
rect -4336 -718 -4278 -706
rect -4218 -130 -4160 -118
rect -4218 -706 -4206 -130
rect -4172 -706 -4160 -130
rect -4218 -718 -4160 -706
rect -4100 -130 -4042 -118
rect -4100 -706 -4088 -130
rect -4054 -706 -4042 -130
rect -4100 -718 -4042 -706
rect -3982 -130 -3924 -118
rect -3982 -706 -3970 -130
rect -3936 -706 -3924 -130
rect -3982 -718 -3924 -706
rect -3864 -130 -3806 -118
rect -3864 -706 -3852 -130
rect -3818 -706 -3806 -130
rect -3864 -718 -3806 -706
rect -3746 -130 -3688 -118
rect -3746 -706 -3734 -130
rect -3700 -706 -3688 -130
rect -3746 -718 -3688 -706
rect -3628 -130 -3570 -118
rect -3628 -706 -3616 -130
rect -3582 -706 -3570 -130
rect -3628 -718 -3570 -706
rect -3510 -130 -3452 -118
rect -3510 -706 -3498 -130
rect -3464 -706 -3452 -130
rect -3510 -718 -3452 -706
rect -3392 -130 -3334 -118
rect -3392 -706 -3380 -130
rect -3346 -706 -3334 -130
rect -3392 -718 -3334 -706
rect -3274 -130 -3216 -118
rect -3274 -706 -3262 -130
rect -3228 -706 -3216 -130
rect -3274 -718 -3216 -706
rect -3156 -130 -3098 -118
rect -3156 -706 -3144 -130
rect -3110 -706 -3098 -130
rect -3156 -718 -3098 -706
rect -3038 -130 -2980 -118
rect -3038 -706 -3026 -130
rect -2992 -706 -2980 -130
rect -3038 -718 -2980 -706
rect -2920 -130 -2862 -118
rect -2920 -706 -2908 -130
rect -2874 -706 -2862 -130
rect -2920 -718 -2862 -706
rect -2802 -130 -2744 -118
rect -2802 -706 -2790 -130
rect -2756 -706 -2744 -130
rect -2802 -718 -2744 -706
rect -2684 -130 -2626 -118
rect -2684 -706 -2672 -130
rect -2638 -706 -2626 -130
rect -2684 -718 -2626 -706
rect -2566 -130 -2508 -118
rect -2566 -706 -2554 -130
rect -2520 -706 -2508 -130
rect -2566 -718 -2508 -706
rect -2448 -130 -2390 -118
rect -2448 -706 -2436 -130
rect -2402 -706 -2390 -130
rect -2448 -718 -2390 -706
rect -2330 -130 -2272 -118
rect -2330 -706 -2318 -130
rect -2284 -706 -2272 -130
rect -2330 -718 -2272 -706
rect -2212 -130 -2154 -118
rect -2212 -706 -2200 -130
rect -2166 -706 -2154 -130
rect -2212 -718 -2154 -706
rect -2094 -130 -2036 -118
rect -2094 -706 -2082 -130
rect -2048 -706 -2036 -130
rect -2094 -718 -2036 -706
rect -1976 -130 -1918 -118
rect -1976 -706 -1964 -130
rect -1930 -706 -1918 -130
rect -1976 -718 -1918 -706
rect -1858 -130 -1800 -118
rect -1858 -706 -1846 -130
rect -1812 -706 -1800 -130
rect -1858 -718 -1800 -706
rect -1740 -130 -1682 -118
rect -1740 -706 -1728 -130
rect -1694 -706 -1682 -130
rect -1740 -718 -1682 -706
rect -1622 -130 -1564 -118
rect -1622 -706 -1610 -130
rect -1576 -706 -1564 -130
rect -1622 -718 -1564 -706
rect -1504 -130 -1446 -118
rect -1504 -706 -1492 -130
rect -1458 -706 -1446 -130
rect -1504 -718 -1446 -706
rect -1386 -130 -1328 -118
rect -1386 -706 -1374 -130
rect -1340 -706 -1328 -130
rect -1386 -718 -1328 -706
rect -1268 -130 -1210 -118
rect -1268 -706 -1256 -130
rect -1222 -706 -1210 -130
rect -1268 -718 -1210 -706
rect -1150 -130 -1092 -118
rect -1150 -706 -1138 -130
rect -1104 -706 -1092 -130
rect -1150 -718 -1092 -706
rect -1032 -130 -974 -118
rect -1032 -706 -1020 -130
rect -986 -706 -974 -130
rect -1032 -718 -974 -706
rect -914 -130 -856 -118
rect -914 -706 -902 -130
rect -868 -706 -856 -130
rect -914 -718 -856 -706
rect -796 -130 -738 -118
rect -796 -706 -784 -130
rect -750 -706 -738 -130
rect -796 -718 -738 -706
rect -678 -130 -620 -118
rect -678 -706 -666 -130
rect -632 -706 -620 -130
rect -678 -718 -620 -706
rect -560 -130 -502 -118
rect -560 -706 -548 -130
rect -514 -706 -502 -130
rect -560 -718 -502 -706
rect -442 -130 -384 -118
rect -442 -706 -430 -130
rect -396 -706 -384 -130
rect -442 -718 -384 -706
rect -324 -130 -266 -118
rect -324 -706 -312 -130
rect -278 -706 -266 -130
rect -324 -718 -266 -706
rect -206 -130 -148 -118
rect -206 -706 -194 -130
rect -160 -706 -148 -130
rect -206 -718 -148 -706
rect -88 -130 -30 -118
rect -88 -706 -76 -130
rect -42 -706 -30 -130
rect -88 -718 -30 -706
rect 30 -130 88 -118
rect 30 -706 42 -130
rect 76 -706 88 -130
rect 30 -718 88 -706
rect 148 -130 206 -118
rect 148 -706 160 -130
rect 194 -706 206 -130
rect 148 -718 206 -706
rect 266 -130 324 -118
rect 266 -706 278 -130
rect 312 -706 324 -130
rect 266 -718 324 -706
rect 384 -130 442 -118
rect 384 -706 396 -130
rect 430 -706 442 -130
rect 384 -718 442 -706
rect 502 -130 560 -118
rect 502 -706 514 -130
rect 548 -706 560 -130
rect 502 -718 560 -706
rect 620 -130 678 -118
rect 620 -706 632 -130
rect 666 -706 678 -130
rect 620 -718 678 -706
rect 738 -130 796 -118
rect 738 -706 750 -130
rect 784 -706 796 -130
rect 738 -718 796 -706
rect 856 -130 914 -118
rect 856 -706 868 -130
rect 902 -706 914 -130
rect 856 -718 914 -706
rect 974 -130 1032 -118
rect 974 -706 986 -130
rect 1020 -706 1032 -130
rect 974 -718 1032 -706
rect 1092 -130 1150 -118
rect 1092 -706 1104 -130
rect 1138 -706 1150 -130
rect 1092 -718 1150 -706
rect 1210 -130 1268 -118
rect 1210 -706 1222 -130
rect 1256 -706 1268 -130
rect 1210 -718 1268 -706
rect 1328 -130 1386 -118
rect 1328 -706 1340 -130
rect 1374 -706 1386 -130
rect 1328 -718 1386 -706
rect 1446 -130 1504 -118
rect 1446 -706 1458 -130
rect 1492 -706 1504 -130
rect 1446 -718 1504 -706
rect 1564 -130 1622 -118
rect 1564 -706 1576 -130
rect 1610 -706 1622 -130
rect 1564 -718 1622 -706
rect 1682 -130 1740 -118
rect 1682 -706 1694 -130
rect 1728 -706 1740 -130
rect 1682 -718 1740 -706
rect 1800 -130 1858 -118
rect 1800 -706 1812 -130
rect 1846 -706 1858 -130
rect 1800 -718 1858 -706
rect 1918 -130 1976 -118
rect 1918 -706 1930 -130
rect 1964 -706 1976 -130
rect 1918 -718 1976 -706
rect 2036 -130 2094 -118
rect 2036 -706 2048 -130
rect 2082 -706 2094 -130
rect 2036 -718 2094 -706
rect 2154 -130 2212 -118
rect 2154 -706 2166 -130
rect 2200 -706 2212 -130
rect 2154 -718 2212 -706
rect 2272 -130 2330 -118
rect 2272 -706 2284 -130
rect 2318 -706 2330 -130
rect 2272 -718 2330 -706
rect 2390 -130 2448 -118
rect 2390 -706 2402 -130
rect 2436 -706 2448 -130
rect 2390 -718 2448 -706
rect 2508 -130 2566 -118
rect 2508 -706 2520 -130
rect 2554 -706 2566 -130
rect 2508 -718 2566 -706
rect 2626 -130 2684 -118
rect 2626 -706 2638 -130
rect 2672 -706 2684 -130
rect 2626 -718 2684 -706
rect 2744 -130 2802 -118
rect 2744 -706 2756 -130
rect 2790 -706 2802 -130
rect 2744 -718 2802 -706
rect 2862 -130 2920 -118
rect 2862 -706 2874 -130
rect 2908 -706 2920 -130
rect 2862 -718 2920 -706
rect 2980 -130 3038 -118
rect 2980 -706 2992 -130
rect 3026 -706 3038 -130
rect 2980 -718 3038 -706
rect 3098 -130 3156 -118
rect 3098 -706 3110 -130
rect 3144 -706 3156 -130
rect 3098 -718 3156 -706
rect 3216 -130 3274 -118
rect 3216 -706 3228 -130
rect 3262 -706 3274 -130
rect 3216 -718 3274 -706
rect 3334 -130 3392 -118
rect 3334 -706 3346 -130
rect 3380 -706 3392 -130
rect 3334 -718 3392 -706
rect 3452 -130 3510 -118
rect 3452 -706 3464 -130
rect 3498 -706 3510 -130
rect 3452 -718 3510 -706
rect 3570 -130 3628 -118
rect 3570 -706 3582 -130
rect 3616 -706 3628 -130
rect 3570 -718 3628 -706
rect 3688 -130 3746 -118
rect 3688 -706 3700 -130
rect 3734 -706 3746 -130
rect 3688 -718 3746 -706
rect 3806 -130 3864 -118
rect 3806 -706 3818 -130
rect 3852 -706 3864 -130
rect 3806 -718 3864 -706
rect 3924 -130 3982 -118
rect 3924 -706 3936 -130
rect 3970 -706 3982 -130
rect 3924 -718 3982 -706
rect 4042 -130 4100 -118
rect 4042 -706 4054 -130
rect 4088 -706 4100 -130
rect 4042 -718 4100 -706
rect 4160 -130 4218 -118
rect 4160 -706 4172 -130
rect 4206 -706 4218 -130
rect 4160 -718 4218 -706
rect 4278 -130 4336 -118
rect 4278 -706 4290 -130
rect 4324 -706 4336 -130
rect 4278 -718 4336 -706
rect 4396 -130 4454 -118
rect 4396 -706 4408 -130
rect 4442 -706 4454 -130
rect 4396 -718 4454 -706
<< pdiffc >>
rect -4442 130 -4408 706
rect -4324 130 -4290 706
rect -4206 130 -4172 706
rect -4088 130 -4054 706
rect -3970 130 -3936 706
rect -3852 130 -3818 706
rect -3734 130 -3700 706
rect -3616 130 -3582 706
rect -3498 130 -3464 706
rect -3380 130 -3346 706
rect -3262 130 -3228 706
rect -3144 130 -3110 706
rect -3026 130 -2992 706
rect -2908 130 -2874 706
rect -2790 130 -2756 706
rect -2672 130 -2638 706
rect -2554 130 -2520 706
rect -2436 130 -2402 706
rect -2318 130 -2284 706
rect -2200 130 -2166 706
rect -2082 130 -2048 706
rect -1964 130 -1930 706
rect -1846 130 -1812 706
rect -1728 130 -1694 706
rect -1610 130 -1576 706
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect 1576 130 1610 706
rect 1694 130 1728 706
rect 1812 130 1846 706
rect 1930 130 1964 706
rect 2048 130 2082 706
rect 2166 130 2200 706
rect 2284 130 2318 706
rect 2402 130 2436 706
rect 2520 130 2554 706
rect 2638 130 2672 706
rect 2756 130 2790 706
rect 2874 130 2908 706
rect 2992 130 3026 706
rect 3110 130 3144 706
rect 3228 130 3262 706
rect 3346 130 3380 706
rect 3464 130 3498 706
rect 3582 130 3616 706
rect 3700 130 3734 706
rect 3818 130 3852 706
rect 3936 130 3970 706
rect 4054 130 4088 706
rect 4172 130 4206 706
rect 4290 130 4324 706
rect 4408 130 4442 706
rect -4442 -706 -4408 -130
rect -4324 -706 -4290 -130
rect -4206 -706 -4172 -130
rect -4088 -706 -4054 -130
rect -3970 -706 -3936 -130
rect -3852 -706 -3818 -130
rect -3734 -706 -3700 -130
rect -3616 -706 -3582 -130
rect -3498 -706 -3464 -130
rect -3380 -706 -3346 -130
rect -3262 -706 -3228 -130
rect -3144 -706 -3110 -130
rect -3026 -706 -2992 -130
rect -2908 -706 -2874 -130
rect -2790 -706 -2756 -130
rect -2672 -706 -2638 -130
rect -2554 -706 -2520 -130
rect -2436 -706 -2402 -130
rect -2318 -706 -2284 -130
rect -2200 -706 -2166 -130
rect -2082 -706 -2048 -130
rect -1964 -706 -1930 -130
rect -1846 -706 -1812 -130
rect -1728 -706 -1694 -130
rect -1610 -706 -1576 -130
rect -1492 -706 -1458 -130
rect -1374 -706 -1340 -130
rect -1256 -706 -1222 -130
rect -1138 -706 -1104 -130
rect -1020 -706 -986 -130
rect -902 -706 -868 -130
rect -784 -706 -750 -130
rect -666 -706 -632 -130
rect -548 -706 -514 -130
rect -430 -706 -396 -130
rect -312 -706 -278 -130
rect -194 -706 -160 -130
rect -76 -706 -42 -130
rect 42 -706 76 -130
rect 160 -706 194 -130
rect 278 -706 312 -130
rect 396 -706 430 -130
rect 514 -706 548 -130
rect 632 -706 666 -130
rect 750 -706 784 -130
rect 868 -706 902 -130
rect 986 -706 1020 -130
rect 1104 -706 1138 -130
rect 1222 -706 1256 -130
rect 1340 -706 1374 -130
rect 1458 -706 1492 -130
rect 1576 -706 1610 -130
rect 1694 -706 1728 -130
rect 1812 -706 1846 -130
rect 1930 -706 1964 -130
rect 2048 -706 2082 -130
rect 2166 -706 2200 -130
rect 2284 -706 2318 -130
rect 2402 -706 2436 -130
rect 2520 -706 2554 -130
rect 2638 -706 2672 -130
rect 2756 -706 2790 -130
rect 2874 -706 2908 -130
rect 2992 -706 3026 -130
rect 3110 -706 3144 -130
rect 3228 -706 3262 -130
rect 3346 -706 3380 -130
rect 3464 -706 3498 -130
rect 3582 -706 3616 -130
rect 3700 -706 3734 -130
rect 3818 -706 3852 -130
rect 3936 -706 3970 -130
rect 4054 -706 4088 -130
rect 4172 -706 4206 -130
rect 4290 -706 4324 -130
rect 4408 -706 4442 -130
<< nsubdiff >>
rect -4556 867 -4460 901
rect 4460 867 4556 901
rect -4556 805 -4522 867
rect 4522 805 4556 867
rect -4556 -867 -4522 -805
rect 4522 -867 4556 -805
rect -4556 -901 -4460 -867
rect 4460 -901 4556 -867
<< nsubdiffcont >>
rect -4460 867 4460 901
rect -4556 -805 -4522 805
rect 4522 -805 4556 805
rect -4460 -901 4460 -867
<< poly >>
rect -4399 799 -4333 815
rect -4399 765 -4383 799
rect -4349 765 -4333 799
rect -4399 749 -4333 765
rect -4281 799 -4215 815
rect -4281 765 -4265 799
rect -4231 765 -4215 799
rect -4281 749 -4215 765
rect -4163 799 -4097 815
rect -4163 765 -4147 799
rect -4113 765 -4097 799
rect -4163 749 -4097 765
rect -4045 799 -3979 815
rect -4045 765 -4029 799
rect -3995 765 -3979 799
rect -4045 749 -3979 765
rect -3927 799 -3861 815
rect -3927 765 -3911 799
rect -3877 765 -3861 799
rect -3927 749 -3861 765
rect -3809 799 -3743 815
rect -3809 765 -3793 799
rect -3759 765 -3743 799
rect -3809 749 -3743 765
rect -3691 799 -3625 815
rect -3691 765 -3675 799
rect -3641 765 -3625 799
rect -3691 749 -3625 765
rect -3573 799 -3507 815
rect -3573 765 -3557 799
rect -3523 765 -3507 799
rect -3573 749 -3507 765
rect -3455 799 -3389 815
rect -3455 765 -3439 799
rect -3405 765 -3389 799
rect -3455 749 -3389 765
rect -3337 799 -3271 815
rect -3337 765 -3321 799
rect -3287 765 -3271 799
rect -3337 749 -3271 765
rect -3219 799 -3153 815
rect -3219 765 -3203 799
rect -3169 765 -3153 799
rect -3219 749 -3153 765
rect -3101 799 -3035 815
rect -3101 765 -3085 799
rect -3051 765 -3035 799
rect -3101 749 -3035 765
rect -2983 799 -2917 815
rect -2983 765 -2967 799
rect -2933 765 -2917 799
rect -2983 749 -2917 765
rect -2865 799 -2799 815
rect -2865 765 -2849 799
rect -2815 765 -2799 799
rect -2865 749 -2799 765
rect -2747 799 -2681 815
rect -2747 765 -2731 799
rect -2697 765 -2681 799
rect -2747 749 -2681 765
rect -2629 799 -2563 815
rect -2629 765 -2613 799
rect -2579 765 -2563 799
rect -2629 749 -2563 765
rect -2511 799 -2445 815
rect -2511 765 -2495 799
rect -2461 765 -2445 799
rect -2511 749 -2445 765
rect -2393 799 -2327 815
rect -2393 765 -2377 799
rect -2343 765 -2327 799
rect -2393 749 -2327 765
rect -2275 799 -2209 815
rect -2275 765 -2259 799
rect -2225 765 -2209 799
rect -2275 749 -2209 765
rect -2157 799 -2091 815
rect -2157 765 -2141 799
rect -2107 765 -2091 799
rect -2157 749 -2091 765
rect -2039 799 -1973 815
rect -2039 765 -2023 799
rect -1989 765 -1973 799
rect -2039 749 -1973 765
rect -1921 799 -1855 815
rect -1921 765 -1905 799
rect -1871 765 -1855 799
rect -1921 749 -1855 765
rect -1803 799 -1737 815
rect -1803 765 -1787 799
rect -1753 765 -1737 799
rect -1803 749 -1737 765
rect -1685 799 -1619 815
rect -1685 765 -1669 799
rect -1635 765 -1619 799
rect -1685 749 -1619 765
rect -1567 799 -1501 815
rect -1567 765 -1551 799
rect -1517 765 -1501 799
rect -1567 749 -1501 765
rect -1449 799 -1383 815
rect -1449 765 -1433 799
rect -1399 765 -1383 799
rect -1449 749 -1383 765
rect -1331 799 -1265 815
rect -1331 765 -1315 799
rect -1281 765 -1265 799
rect -1331 749 -1265 765
rect -1213 799 -1147 815
rect -1213 765 -1197 799
rect -1163 765 -1147 799
rect -1213 749 -1147 765
rect -1095 799 -1029 815
rect -1095 765 -1079 799
rect -1045 765 -1029 799
rect -1095 749 -1029 765
rect -977 799 -911 815
rect -977 765 -961 799
rect -927 765 -911 799
rect -977 749 -911 765
rect -859 799 -793 815
rect -859 765 -843 799
rect -809 765 -793 799
rect -859 749 -793 765
rect -741 799 -675 815
rect -741 765 -725 799
rect -691 765 -675 799
rect -741 749 -675 765
rect -623 799 -557 815
rect -623 765 -607 799
rect -573 765 -557 799
rect -623 749 -557 765
rect -505 799 -439 815
rect -505 765 -489 799
rect -455 765 -439 799
rect -505 749 -439 765
rect -387 799 -321 815
rect -387 765 -371 799
rect -337 765 -321 799
rect -387 749 -321 765
rect -269 799 -203 815
rect -269 765 -253 799
rect -219 765 -203 799
rect -269 749 -203 765
rect -151 799 -85 815
rect -151 765 -135 799
rect -101 765 -85 799
rect -151 749 -85 765
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect 85 799 151 815
rect 85 765 101 799
rect 135 765 151 799
rect 85 749 151 765
rect 203 799 269 815
rect 203 765 219 799
rect 253 765 269 799
rect 203 749 269 765
rect 321 799 387 815
rect 321 765 337 799
rect 371 765 387 799
rect 321 749 387 765
rect 439 799 505 815
rect 439 765 455 799
rect 489 765 505 799
rect 439 749 505 765
rect 557 799 623 815
rect 557 765 573 799
rect 607 765 623 799
rect 557 749 623 765
rect 675 799 741 815
rect 675 765 691 799
rect 725 765 741 799
rect 675 749 741 765
rect 793 799 859 815
rect 793 765 809 799
rect 843 765 859 799
rect 793 749 859 765
rect 911 799 977 815
rect 911 765 927 799
rect 961 765 977 799
rect 911 749 977 765
rect 1029 799 1095 815
rect 1029 765 1045 799
rect 1079 765 1095 799
rect 1029 749 1095 765
rect 1147 799 1213 815
rect 1147 765 1163 799
rect 1197 765 1213 799
rect 1147 749 1213 765
rect 1265 799 1331 815
rect 1265 765 1281 799
rect 1315 765 1331 799
rect 1265 749 1331 765
rect 1383 799 1449 815
rect 1383 765 1399 799
rect 1433 765 1449 799
rect 1383 749 1449 765
rect 1501 799 1567 815
rect 1501 765 1517 799
rect 1551 765 1567 799
rect 1501 749 1567 765
rect 1619 799 1685 815
rect 1619 765 1635 799
rect 1669 765 1685 799
rect 1619 749 1685 765
rect 1737 799 1803 815
rect 1737 765 1753 799
rect 1787 765 1803 799
rect 1737 749 1803 765
rect 1855 799 1921 815
rect 1855 765 1871 799
rect 1905 765 1921 799
rect 1855 749 1921 765
rect 1973 799 2039 815
rect 1973 765 1989 799
rect 2023 765 2039 799
rect 1973 749 2039 765
rect 2091 799 2157 815
rect 2091 765 2107 799
rect 2141 765 2157 799
rect 2091 749 2157 765
rect 2209 799 2275 815
rect 2209 765 2225 799
rect 2259 765 2275 799
rect 2209 749 2275 765
rect 2327 799 2393 815
rect 2327 765 2343 799
rect 2377 765 2393 799
rect 2327 749 2393 765
rect 2445 799 2511 815
rect 2445 765 2461 799
rect 2495 765 2511 799
rect 2445 749 2511 765
rect 2563 799 2629 815
rect 2563 765 2579 799
rect 2613 765 2629 799
rect 2563 749 2629 765
rect 2681 799 2747 815
rect 2681 765 2697 799
rect 2731 765 2747 799
rect 2681 749 2747 765
rect 2799 799 2865 815
rect 2799 765 2815 799
rect 2849 765 2865 799
rect 2799 749 2865 765
rect 2917 799 2983 815
rect 2917 765 2933 799
rect 2967 765 2983 799
rect 2917 749 2983 765
rect 3035 799 3101 815
rect 3035 765 3051 799
rect 3085 765 3101 799
rect 3035 749 3101 765
rect 3153 799 3219 815
rect 3153 765 3169 799
rect 3203 765 3219 799
rect 3153 749 3219 765
rect 3271 799 3337 815
rect 3271 765 3287 799
rect 3321 765 3337 799
rect 3271 749 3337 765
rect 3389 799 3455 815
rect 3389 765 3405 799
rect 3439 765 3455 799
rect 3389 749 3455 765
rect 3507 799 3573 815
rect 3507 765 3523 799
rect 3557 765 3573 799
rect 3507 749 3573 765
rect 3625 799 3691 815
rect 3625 765 3641 799
rect 3675 765 3691 799
rect 3625 749 3691 765
rect 3743 799 3809 815
rect 3743 765 3759 799
rect 3793 765 3809 799
rect 3743 749 3809 765
rect 3861 799 3927 815
rect 3861 765 3877 799
rect 3911 765 3927 799
rect 3861 749 3927 765
rect 3979 799 4045 815
rect 3979 765 3995 799
rect 4029 765 4045 799
rect 3979 749 4045 765
rect 4097 799 4163 815
rect 4097 765 4113 799
rect 4147 765 4163 799
rect 4097 749 4163 765
rect 4215 799 4281 815
rect 4215 765 4231 799
rect 4265 765 4281 799
rect 4215 749 4281 765
rect 4333 799 4399 815
rect 4333 765 4349 799
rect 4383 765 4399 799
rect 4333 749 4399 765
rect -4396 718 -4336 749
rect -4278 718 -4218 749
rect -4160 718 -4100 749
rect -4042 718 -3982 749
rect -3924 718 -3864 749
rect -3806 718 -3746 749
rect -3688 718 -3628 749
rect -3570 718 -3510 749
rect -3452 718 -3392 749
rect -3334 718 -3274 749
rect -3216 718 -3156 749
rect -3098 718 -3038 749
rect -2980 718 -2920 749
rect -2862 718 -2802 749
rect -2744 718 -2684 749
rect -2626 718 -2566 749
rect -2508 718 -2448 749
rect -2390 718 -2330 749
rect -2272 718 -2212 749
rect -2154 718 -2094 749
rect -2036 718 -1976 749
rect -1918 718 -1858 749
rect -1800 718 -1740 749
rect -1682 718 -1622 749
rect -1564 718 -1504 749
rect -1446 718 -1386 749
rect -1328 718 -1268 749
rect -1210 718 -1150 749
rect -1092 718 -1032 749
rect -974 718 -914 749
rect -856 718 -796 749
rect -738 718 -678 749
rect -620 718 -560 749
rect -502 718 -442 749
rect -384 718 -324 749
rect -266 718 -206 749
rect -148 718 -88 749
rect -30 718 30 749
rect 88 718 148 749
rect 206 718 266 749
rect 324 718 384 749
rect 442 718 502 749
rect 560 718 620 749
rect 678 718 738 749
rect 796 718 856 749
rect 914 718 974 749
rect 1032 718 1092 749
rect 1150 718 1210 749
rect 1268 718 1328 749
rect 1386 718 1446 749
rect 1504 718 1564 749
rect 1622 718 1682 749
rect 1740 718 1800 749
rect 1858 718 1918 749
rect 1976 718 2036 749
rect 2094 718 2154 749
rect 2212 718 2272 749
rect 2330 718 2390 749
rect 2448 718 2508 749
rect 2566 718 2626 749
rect 2684 718 2744 749
rect 2802 718 2862 749
rect 2920 718 2980 749
rect 3038 718 3098 749
rect 3156 718 3216 749
rect 3274 718 3334 749
rect 3392 718 3452 749
rect 3510 718 3570 749
rect 3628 718 3688 749
rect 3746 718 3806 749
rect 3864 718 3924 749
rect 3982 718 4042 749
rect 4100 718 4160 749
rect 4218 718 4278 749
rect 4336 718 4396 749
rect -4396 87 -4336 118
rect -4278 87 -4218 118
rect -4160 87 -4100 118
rect -4042 87 -3982 118
rect -3924 87 -3864 118
rect -3806 87 -3746 118
rect -3688 87 -3628 118
rect -3570 87 -3510 118
rect -3452 87 -3392 118
rect -3334 87 -3274 118
rect -3216 87 -3156 118
rect -3098 87 -3038 118
rect -2980 87 -2920 118
rect -2862 87 -2802 118
rect -2744 87 -2684 118
rect -2626 87 -2566 118
rect -2508 87 -2448 118
rect -2390 87 -2330 118
rect -2272 87 -2212 118
rect -2154 87 -2094 118
rect -2036 87 -1976 118
rect -1918 87 -1858 118
rect -1800 87 -1740 118
rect -1682 87 -1622 118
rect -1564 87 -1504 118
rect -1446 87 -1386 118
rect -1328 87 -1268 118
rect -1210 87 -1150 118
rect -1092 87 -1032 118
rect -974 87 -914 118
rect -856 87 -796 118
rect -738 87 -678 118
rect -620 87 -560 118
rect -502 87 -442 118
rect -384 87 -324 118
rect -266 87 -206 118
rect -148 87 -88 118
rect -30 87 30 118
rect 88 87 148 118
rect 206 87 266 118
rect 324 87 384 118
rect 442 87 502 118
rect 560 87 620 118
rect 678 87 738 118
rect 796 87 856 118
rect 914 87 974 118
rect 1032 87 1092 118
rect 1150 87 1210 118
rect 1268 87 1328 118
rect 1386 87 1446 118
rect 1504 87 1564 118
rect 1622 87 1682 118
rect 1740 87 1800 118
rect 1858 87 1918 118
rect 1976 87 2036 118
rect 2094 87 2154 118
rect 2212 87 2272 118
rect 2330 87 2390 118
rect 2448 87 2508 118
rect 2566 87 2626 118
rect 2684 87 2744 118
rect 2802 87 2862 118
rect 2920 87 2980 118
rect 3038 87 3098 118
rect 3156 87 3216 118
rect 3274 87 3334 118
rect 3392 87 3452 118
rect 3510 87 3570 118
rect 3628 87 3688 118
rect 3746 87 3806 118
rect 3864 87 3924 118
rect 3982 87 4042 118
rect 4100 87 4160 118
rect 4218 87 4278 118
rect 4336 87 4396 118
rect -4399 71 -4333 87
rect -4399 37 -4383 71
rect -4349 37 -4333 71
rect -4399 21 -4333 37
rect -4281 71 -4215 87
rect -4281 37 -4265 71
rect -4231 37 -4215 71
rect -4281 21 -4215 37
rect -4163 71 -4097 87
rect -4163 37 -4147 71
rect -4113 37 -4097 71
rect -4163 21 -4097 37
rect -4045 71 -3979 87
rect -4045 37 -4029 71
rect -3995 37 -3979 71
rect -4045 21 -3979 37
rect -3927 71 -3861 87
rect -3927 37 -3911 71
rect -3877 37 -3861 71
rect -3927 21 -3861 37
rect -3809 71 -3743 87
rect -3809 37 -3793 71
rect -3759 37 -3743 71
rect -3809 21 -3743 37
rect -3691 71 -3625 87
rect -3691 37 -3675 71
rect -3641 37 -3625 71
rect -3691 21 -3625 37
rect -3573 71 -3507 87
rect -3573 37 -3557 71
rect -3523 37 -3507 71
rect -3573 21 -3507 37
rect -3455 71 -3389 87
rect -3455 37 -3439 71
rect -3405 37 -3389 71
rect -3455 21 -3389 37
rect -3337 71 -3271 87
rect -3337 37 -3321 71
rect -3287 37 -3271 71
rect -3337 21 -3271 37
rect -3219 71 -3153 87
rect -3219 37 -3203 71
rect -3169 37 -3153 71
rect -3219 21 -3153 37
rect -3101 71 -3035 87
rect -3101 37 -3085 71
rect -3051 37 -3035 71
rect -3101 21 -3035 37
rect -2983 71 -2917 87
rect -2983 37 -2967 71
rect -2933 37 -2917 71
rect -2983 21 -2917 37
rect -2865 71 -2799 87
rect -2865 37 -2849 71
rect -2815 37 -2799 71
rect -2865 21 -2799 37
rect -2747 71 -2681 87
rect -2747 37 -2731 71
rect -2697 37 -2681 71
rect -2747 21 -2681 37
rect -2629 71 -2563 87
rect -2629 37 -2613 71
rect -2579 37 -2563 71
rect -2629 21 -2563 37
rect -2511 71 -2445 87
rect -2511 37 -2495 71
rect -2461 37 -2445 71
rect -2511 21 -2445 37
rect -2393 71 -2327 87
rect -2393 37 -2377 71
rect -2343 37 -2327 71
rect -2393 21 -2327 37
rect -2275 71 -2209 87
rect -2275 37 -2259 71
rect -2225 37 -2209 71
rect -2275 21 -2209 37
rect -2157 71 -2091 87
rect -2157 37 -2141 71
rect -2107 37 -2091 71
rect -2157 21 -2091 37
rect -2039 71 -1973 87
rect -2039 37 -2023 71
rect -1989 37 -1973 71
rect -2039 21 -1973 37
rect -1921 71 -1855 87
rect -1921 37 -1905 71
rect -1871 37 -1855 71
rect -1921 21 -1855 37
rect -1803 71 -1737 87
rect -1803 37 -1787 71
rect -1753 37 -1737 71
rect -1803 21 -1737 37
rect -1685 71 -1619 87
rect -1685 37 -1669 71
rect -1635 37 -1619 71
rect -1685 21 -1619 37
rect -1567 71 -1501 87
rect -1567 37 -1551 71
rect -1517 37 -1501 71
rect -1567 21 -1501 37
rect -1449 71 -1383 87
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1449 21 -1383 37
rect -1331 71 -1265 87
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1331 21 -1265 37
rect -1213 71 -1147 87
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1213 21 -1147 37
rect -1095 71 -1029 87
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -1095 21 -1029 37
rect -977 71 -911 87
rect -977 37 -961 71
rect -927 37 -911 71
rect -977 21 -911 37
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect 911 71 977 87
rect 911 37 927 71
rect 961 37 977 71
rect 911 21 977 37
rect 1029 71 1095 87
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1029 21 1095 37
rect 1147 71 1213 87
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1147 21 1213 37
rect 1265 71 1331 87
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1265 21 1331 37
rect 1383 71 1449 87
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1383 21 1449 37
rect 1501 71 1567 87
rect 1501 37 1517 71
rect 1551 37 1567 71
rect 1501 21 1567 37
rect 1619 71 1685 87
rect 1619 37 1635 71
rect 1669 37 1685 71
rect 1619 21 1685 37
rect 1737 71 1803 87
rect 1737 37 1753 71
rect 1787 37 1803 71
rect 1737 21 1803 37
rect 1855 71 1921 87
rect 1855 37 1871 71
rect 1905 37 1921 71
rect 1855 21 1921 37
rect 1973 71 2039 87
rect 1973 37 1989 71
rect 2023 37 2039 71
rect 1973 21 2039 37
rect 2091 71 2157 87
rect 2091 37 2107 71
rect 2141 37 2157 71
rect 2091 21 2157 37
rect 2209 71 2275 87
rect 2209 37 2225 71
rect 2259 37 2275 71
rect 2209 21 2275 37
rect 2327 71 2393 87
rect 2327 37 2343 71
rect 2377 37 2393 71
rect 2327 21 2393 37
rect 2445 71 2511 87
rect 2445 37 2461 71
rect 2495 37 2511 71
rect 2445 21 2511 37
rect 2563 71 2629 87
rect 2563 37 2579 71
rect 2613 37 2629 71
rect 2563 21 2629 37
rect 2681 71 2747 87
rect 2681 37 2697 71
rect 2731 37 2747 71
rect 2681 21 2747 37
rect 2799 71 2865 87
rect 2799 37 2815 71
rect 2849 37 2865 71
rect 2799 21 2865 37
rect 2917 71 2983 87
rect 2917 37 2933 71
rect 2967 37 2983 71
rect 2917 21 2983 37
rect 3035 71 3101 87
rect 3035 37 3051 71
rect 3085 37 3101 71
rect 3035 21 3101 37
rect 3153 71 3219 87
rect 3153 37 3169 71
rect 3203 37 3219 71
rect 3153 21 3219 37
rect 3271 71 3337 87
rect 3271 37 3287 71
rect 3321 37 3337 71
rect 3271 21 3337 37
rect 3389 71 3455 87
rect 3389 37 3405 71
rect 3439 37 3455 71
rect 3389 21 3455 37
rect 3507 71 3573 87
rect 3507 37 3523 71
rect 3557 37 3573 71
rect 3507 21 3573 37
rect 3625 71 3691 87
rect 3625 37 3641 71
rect 3675 37 3691 71
rect 3625 21 3691 37
rect 3743 71 3809 87
rect 3743 37 3759 71
rect 3793 37 3809 71
rect 3743 21 3809 37
rect 3861 71 3927 87
rect 3861 37 3877 71
rect 3911 37 3927 71
rect 3861 21 3927 37
rect 3979 71 4045 87
rect 3979 37 3995 71
rect 4029 37 4045 71
rect 3979 21 4045 37
rect 4097 71 4163 87
rect 4097 37 4113 71
rect 4147 37 4163 71
rect 4097 21 4163 37
rect 4215 71 4281 87
rect 4215 37 4231 71
rect 4265 37 4281 71
rect 4215 21 4281 37
rect 4333 71 4399 87
rect 4333 37 4349 71
rect 4383 37 4399 71
rect 4333 21 4399 37
rect -4399 -37 -4333 -21
rect -4399 -71 -4383 -37
rect -4349 -71 -4333 -37
rect -4399 -87 -4333 -71
rect -4281 -37 -4215 -21
rect -4281 -71 -4265 -37
rect -4231 -71 -4215 -37
rect -4281 -87 -4215 -71
rect -4163 -37 -4097 -21
rect -4163 -71 -4147 -37
rect -4113 -71 -4097 -37
rect -4163 -87 -4097 -71
rect -4045 -37 -3979 -21
rect -4045 -71 -4029 -37
rect -3995 -71 -3979 -37
rect -4045 -87 -3979 -71
rect -3927 -37 -3861 -21
rect -3927 -71 -3911 -37
rect -3877 -71 -3861 -37
rect -3927 -87 -3861 -71
rect -3809 -37 -3743 -21
rect -3809 -71 -3793 -37
rect -3759 -71 -3743 -37
rect -3809 -87 -3743 -71
rect -3691 -37 -3625 -21
rect -3691 -71 -3675 -37
rect -3641 -71 -3625 -37
rect -3691 -87 -3625 -71
rect -3573 -37 -3507 -21
rect -3573 -71 -3557 -37
rect -3523 -71 -3507 -37
rect -3573 -87 -3507 -71
rect -3455 -37 -3389 -21
rect -3455 -71 -3439 -37
rect -3405 -71 -3389 -37
rect -3455 -87 -3389 -71
rect -3337 -37 -3271 -21
rect -3337 -71 -3321 -37
rect -3287 -71 -3271 -37
rect -3337 -87 -3271 -71
rect -3219 -37 -3153 -21
rect -3219 -71 -3203 -37
rect -3169 -71 -3153 -37
rect -3219 -87 -3153 -71
rect -3101 -37 -3035 -21
rect -3101 -71 -3085 -37
rect -3051 -71 -3035 -37
rect -3101 -87 -3035 -71
rect -2983 -37 -2917 -21
rect -2983 -71 -2967 -37
rect -2933 -71 -2917 -37
rect -2983 -87 -2917 -71
rect -2865 -37 -2799 -21
rect -2865 -71 -2849 -37
rect -2815 -71 -2799 -37
rect -2865 -87 -2799 -71
rect -2747 -37 -2681 -21
rect -2747 -71 -2731 -37
rect -2697 -71 -2681 -37
rect -2747 -87 -2681 -71
rect -2629 -37 -2563 -21
rect -2629 -71 -2613 -37
rect -2579 -71 -2563 -37
rect -2629 -87 -2563 -71
rect -2511 -37 -2445 -21
rect -2511 -71 -2495 -37
rect -2461 -71 -2445 -37
rect -2511 -87 -2445 -71
rect -2393 -37 -2327 -21
rect -2393 -71 -2377 -37
rect -2343 -71 -2327 -37
rect -2393 -87 -2327 -71
rect -2275 -37 -2209 -21
rect -2275 -71 -2259 -37
rect -2225 -71 -2209 -37
rect -2275 -87 -2209 -71
rect -2157 -37 -2091 -21
rect -2157 -71 -2141 -37
rect -2107 -71 -2091 -37
rect -2157 -87 -2091 -71
rect -2039 -37 -1973 -21
rect -2039 -71 -2023 -37
rect -1989 -71 -1973 -37
rect -2039 -87 -1973 -71
rect -1921 -37 -1855 -21
rect -1921 -71 -1905 -37
rect -1871 -71 -1855 -37
rect -1921 -87 -1855 -71
rect -1803 -37 -1737 -21
rect -1803 -71 -1787 -37
rect -1753 -71 -1737 -37
rect -1803 -87 -1737 -71
rect -1685 -37 -1619 -21
rect -1685 -71 -1669 -37
rect -1635 -71 -1619 -37
rect -1685 -87 -1619 -71
rect -1567 -37 -1501 -21
rect -1567 -71 -1551 -37
rect -1517 -71 -1501 -37
rect -1567 -87 -1501 -71
rect -1449 -37 -1383 -21
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1449 -87 -1383 -71
rect -1331 -37 -1265 -21
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1331 -87 -1265 -71
rect -1213 -37 -1147 -21
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1213 -87 -1147 -71
rect -1095 -37 -1029 -21
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -1095 -87 -1029 -71
rect -977 -37 -911 -21
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -977 -87 -911 -71
rect -859 -37 -793 -21
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -859 -87 -793 -71
rect -741 -37 -675 -21
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -741 -87 -675 -71
rect -623 -37 -557 -21
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -623 -87 -557 -71
rect -505 -37 -439 -21
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -505 -87 -439 -71
rect -387 -37 -321 -21
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -387 -87 -321 -71
rect -269 -37 -203 -21
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -269 -87 -203 -71
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect 203 -37 269 -21
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 203 -87 269 -71
rect 321 -37 387 -21
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 321 -87 387 -71
rect 439 -37 505 -21
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 439 -87 505 -71
rect 557 -37 623 -21
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 557 -87 623 -71
rect 675 -37 741 -21
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 675 -87 741 -71
rect 793 -37 859 -21
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 793 -87 859 -71
rect 911 -37 977 -21
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 911 -87 977 -71
rect 1029 -37 1095 -21
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1029 -87 1095 -71
rect 1147 -37 1213 -21
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1147 -87 1213 -71
rect 1265 -37 1331 -21
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1265 -87 1331 -71
rect 1383 -37 1449 -21
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect 1383 -87 1449 -71
rect 1501 -37 1567 -21
rect 1501 -71 1517 -37
rect 1551 -71 1567 -37
rect 1501 -87 1567 -71
rect 1619 -37 1685 -21
rect 1619 -71 1635 -37
rect 1669 -71 1685 -37
rect 1619 -87 1685 -71
rect 1737 -37 1803 -21
rect 1737 -71 1753 -37
rect 1787 -71 1803 -37
rect 1737 -87 1803 -71
rect 1855 -37 1921 -21
rect 1855 -71 1871 -37
rect 1905 -71 1921 -37
rect 1855 -87 1921 -71
rect 1973 -37 2039 -21
rect 1973 -71 1989 -37
rect 2023 -71 2039 -37
rect 1973 -87 2039 -71
rect 2091 -37 2157 -21
rect 2091 -71 2107 -37
rect 2141 -71 2157 -37
rect 2091 -87 2157 -71
rect 2209 -37 2275 -21
rect 2209 -71 2225 -37
rect 2259 -71 2275 -37
rect 2209 -87 2275 -71
rect 2327 -37 2393 -21
rect 2327 -71 2343 -37
rect 2377 -71 2393 -37
rect 2327 -87 2393 -71
rect 2445 -37 2511 -21
rect 2445 -71 2461 -37
rect 2495 -71 2511 -37
rect 2445 -87 2511 -71
rect 2563 -37 2629 -21
rect 2563 -71 2579 -37
rect 2613 -71 2629 -37
rect 2563 -87 2629 -71
rect 2681 -37 2747 -21
rect 2681 -71 2697 -37
rect 2731 -71 2747 -37
rect 2681 -87 2747 -71
rect 2799 -37 2865 -21
rect 2799 -71 2815 -37
rect 2849 -71 2865 -37
rect 2799 -87 2865 -71
rect 2917 -37 2983 -21
rect 2917 -71 2933 -37
rect 2967 -71 2983 -37
rect 2917 -87 2983 -71
rect 3035 -37 3101 -21
rect 3035 -71 3051 -37
rect 3085 -71 3101 -37
rect 3035 -87 3101 -71
rect 3153 -37 3219 -21
rect 3153 -71 3169 -37
rect 3203 -71 3219 -37
rect 3153 -87 3219 -71
rect 3271 -37 3337 -21
rect 3271 -71 3287 -37
rect 3321 -71 3337 -37
rect 3271 -87 3337 -71
rect 3389 -37 3455 -21
rect 3389 -71 3405 -37
rect 3439 -71 3455 -37
rect 3389 -87 3455 -71
rect 3507 -37 3573 -21
rect 3507 -71 3523 -37
rect 3557 -71 3573 -37
rect 3507 -87 3573 -71
rect 3625 -37 3691 -21
rect 3625 -71 3641 -37
rect 3675 -71 3691 -37
rect 3625 -87 3691 -71
rect 3743 -37 3809 -21
rect 3743 -71 3759 -37
rect 3793 -71 3809 -37
rect 3743 -87 3809 -71
rect 3861 -37 3927 -21
rect 3861 -71 3877 -37
rect 3911 -71 3927 -37
rect 3861 -87 3927 -71
rect 3979 -37 4045 -21
rect 3979 -71 3995 -37
rect 4029 -71 4045 -37
rect 3979 -87 4045 -71
rect 4097 -37 4163 -21
rect 4097 -71 4113 -37
rect 4147 -71 4163 -37
rect 4097 -87 4163 -71
rect 4215 -37 4281 -21
rect 4215 -71 4231 -37
rect 4265 -71 4281 -37
rect 4215 -87 4281 -71
rect 4333 -37 4399 -21
rect 4333 -71 4349 -37
rect 4383 -71 4399 -37
rect 4333 -87 4399 -71
rect -4396 -118 -4336 -87
rect -4278 -118 -4218 -87
rect -4160 -118 -4100 -87
rect -4042 -118 -3982 -87
rect -3924 -118 -3864 -87
rect -3806 -118 -3746 -87
rect -3688 -118 -3628 -87
rect -3570 -118 -3510 -87
rect -3452 -118 -3392 -87
rect -3334 -118 -3274 -87
rect -3216 -118 -3156 -87
rect -3098 -118 -3038 -87
rect -2980 -118 -2920 -87
rect -2862 -118 -2802 -87
rect -2744 -118 -2684 -87
rect -2626 -118 -2566 -87
rect -2508 -118 -2448 -87
rect -2390 -118 -2330 -87
rect -2272 -118 -2212 -87
rect -2154 -118 -2094 -87
rect -2036 -118 -1976 -87
rect -1918 -118 -1858 -87
rect -1800 -118 -1740 -87
rect -1682 -118 -1622 -87
rect -1564 -118 -1504 -87
rect -1446 -118 -1386 -87
rect -1328 -118 -1268 -87
rect -1210 -118 -1150 -87
rect -1092 -118 -1032 -87
rect -974 -118 -914 -87
rect -856 -118 -796 -87
rect -738 -118 -678 -87
rect -620 -118 -560 -87
rect -502 -118 -442 -87
rect -384 -118 -324 -87
rect -266 -118 -206 -87
rect -148 -118 -88 -87
rect -30 -118 30 -87
rect 88 -118 148 -87
rect 206 -118 266 -87
rect 324 -118 384 -87
rect 442 -118 502 -87
rect 560 -118 620 -87
rect 678 -118 738 -87
rect 796 -118 856 -87
rect 914 -118 974 -87
rect 1032 -118 1092 -87
rect 1150 -118 1210 -87
rect 1268 -118 1328 -87
rect 1386 -118 1446 -87
rect 1504 -118 1564 -87
rect 1622 -118 1682 -87
rect 1740 -118 1800 -87
rect 1858 -118 1918 -87
rect 1976 -118 2036 -87
rect 2094 -118 2154 -87
rect 2212 -118 2272 -87
rect 2330 -118 2390 -87
rect 2448 -118 2508 -87
rect 2566 -118 2626 -87
rect 2684 -118 2744 -87
rect 2802 -118 2862 -87
rect 2920 -118 2980 -87
rect 3038 -118 3098 -87
rect 3156 -118 3216 -87
rect 3274 -118 3334 -87
rect 3392 -118 3452 -87
rect 3510 -118 3570 -87
rect 3628 -118 3688 -87
rect 3746 -118 3806 -87
rect 3864 -118 3924 -87
rect 3982 -118 4042 -87
rect 4100 -118 4160 -87
rect 4218 -118 4278 -87
rect 4336 -118 4396 -87
rect -4396 -749 -4336 -718
rect -4278 -749 -4218 -718
rect -4160 -749 -4100 -718
rect -4042 -749 -3982 -718
rect -3924 -749 -3864 -718
rect -3806 -749 -3746 -718
rect -3688 -749 -3628 -718
rect -3570 -749 -3510 -718
rect -3452 -749 -3392 -718
rect -3334 -749 -3274 -718
rect -3216 -749 -3156 -718
rect -3098 -749 -3038 -718
rect -2980 -749 -2920 -718
rect -2862 -749 -2802 -718
rect -2744 -749 -2684 -718
rect -2626 -749 -2566 -718
rect -2508 -749 -2448 -718
rect -2390 -749 -2330 -718
rect -2272 -749 -2212 -718
rect -2154 -749 -2094 -718
rect -2036 -749 -1976 -718
rect -1918 -749 -1858 -718
rect -1800 -749 -1740 -718
rect -1682 -749 -1622 -718
rect -1564 -749 -1504 -718
rect -1446 -749 -1386 -718
rect -1328 -749 -1268 -718
rect -1210 -749 -1150 -718
rect -1092 -749 -1032 -718
rect -974 -749 -914 -718
rect -856 -749 -796 -718
rect -738 -749 -678 -718
rect -620 -749 -560 -718
rect -502 -749 -442 -718
rect -384 -749 -324 -718
rect -266 -749 -206 -718
rect -148 -749 -88 -718
rect -30 -749 30 -718
rect 88 -749 148 -718
rect 206 -749 266 -718
rect 324 -749 384 -718
rect 442 -749 502 -718
rect 560 -749 620 -718
rect 678 -749 738 -718
rect 796 -749 856 -718
rect 914 -749 974 -718
rect 1032 -749 1092 -718
rect 1150 -749 1210 -718
rect 1268 -749 1328 -718
rect 1386 -749 1446 -718
rect 1504 -749 1564 -718
rect 1622 -749 1682 -718
rect 1740 -749 1800 -718
rect 1858 -749 1918 -718
rect 1976 -749 2036 -718
rect 2094 -749 2154 -718
rect 2212 -749 2272 -718
rect 2330 -749 2390 -718
rect 2448 -749 2508 -718
rect 2566 -749 2626 -718
rect 2684 -749 2744 -718
rect 2802 -749 2862 -718
rect 2920 -749 2980 -718
rect 3038 -749 3098 -718
rect 3156 -749 3216 -718
rect 3274 -749 3334 -718
rect 3392 -749 3452 -718
rect 3510 -749 3570 -718
rect 3628 -749 3688 -718
rect 3746 -749 3806 -718
rect 3864 -749 3924 -718
rect 3982 -749 4042 -718
rect 4100 -749 4160 -718
rect 4218 -749 4278 -718
rect 4336 -749 4396 -718
rect -4399 -765 -4333 -749
rect -4399 -799 -4383 -765
rect -4349 -799 -4333 -765
rect -4399 -815 -4333 -799
rect -4281 -765 -4215 -749
rect -4281 -799 -4265 -765
rect -4231 -799 -4215 -765
rect -4281 -815 -4215 -799
rect -4163 -765 -4097 -749
rect -4163 -799 -4147 -765
rect -4113 -799 -4097 -765
rect -4163 -815 -4097 -799
rect -4045 -765 -3979 -749
rect -4045 -799 -4029 -765
rect -3995 -799 -3979 -765
rect -4045 -815 -3979 -799
rect -3927 -765 -3861 -749
rect -3927 -799 -3911 -765
rect -3877 -799 -3861 -765
rect -3927 -815 -3861 -799
rect -3809 -765 -3743 -749
rect -3809 -799 -3793 -765
rect -3759 -799 -3743 -765
rect -3809 -815 -3743 -799
rect -3691 -765 -3625 -749
rect -3691 -799 -3675 -765
rect -3641 -799 -3625 -765
rect -3691 -815 -3625 -799
rect -3573 -765 -3507 -749
rect -3573 -799 -3557 -765
rect -3523 -799 -3507 -765
rect -3573 -815 -3507 -799
rect -3455 -765 -3389 -749
rect -3455 -799 -3439 -765
rect -3405 -799 -3389 -765
rect -3455 -815 -3389 -799
rect -3337 -765 -3271 -749
rect -3337 -799 -3321 -765
rect -3287 -799 -3271 -765
rect -3337 -815 -3271 -799
rect -3219 -765 -3153 -749
rect -3219 -799 -3203 -765
rect -3169 -799 -3153 -765
rect -3219 -815 -3153 -799
rect -3101 -765 -3035 -749
rect -3101 -799 -3085 -765
rect -3051 -799 -3035 -765
rect -3101 -815 -3035 -799
rect -2983 -765 -2917 -749
rect -2983 -799 -2967 -765
rect -2933 -799 -2917 -765
rect -2983 -815 -2917 -799
rect -2865 -765 -2799 -749
rect -2865 -799 -2849 -765
rect -2815 -799 -2799 -765
rect -2865 -815 -2799 -799
rect -2747 -765 -2681 -749
rect -2747 -799 -2731 -765
rect -2697 -799 -2681 -765
rect -2747 -815 -2681 -799
rect -2629 -765 -2563 -749
rect -2629 -799 -2613 -765
rect -2579 -799 -2563 -765
rect -2629 -815 -2563 -799
rect -2511 -765 -2445 -749
rect -2511 -799 -2495 -765
rect -2461 -799 -2445 -765
rect -2511 -815 -2445 -799
rect -2393 -765 -2327 -749
rect -2393 -799 -2377 -765
rect -2343 -799 -2327 -765
rect -2393 -815 -2327 -799
rect -2275 -765 -2209 -749
rect -2275 -799 -2259 -765
rect -2225 -799 -2209 -765
rect -2275 -815 -2209 -799
rect -2157 -765 -2091 -749
rect -2157 -799 -2141 -765
rect -2107 -799 -2091 -765
rect -2157 -815 -2091 -799
rect -2039 -765 -1973 -749
rect -2039 -799 -2023 -765
rect -1989 -799 -1973 -765
rect -2039 -815 -1973 -799
rect -1921 -765 -1855 -749
rect -1921 -799 -1905 -765
rect -1871 -799 -1855 -765
rect -1921 -815 -1855 -799
rect -1803 -765 -1737 -749
rect -1803 -799 -1787 -765
rect -1753 -799 -1737 -765
rect -1803 -815 -1737 -799
rect -1685 -765 -1619 -749
rect -1685 -799 -1669 -765
rect -1635 -799 -1619 -765
rect -1685 -815 -1619 -799
rect -1567 -765 -1501 -749
rect -1567 -799 -1551 -765
rect -1517 -799 -1501 -765
rect -1567 -815 -1501 -799
rect -1449 -765 -1383 -749
rect -1449 -799 -1433 -765
rect -1399 -799 -1383 -765
rect -1449 -815 -1383 -799
rect -1331 -765 -1265 -749
rect -1331 -799 -1315 -765
rect -1281 -799 -1265 -765
rect -1331 -815 -1265 -799
rect -1213 -765 -1147 -749
rect -1213 -799 -1197 -765
rect -1163 -799 -1147 -765
rect -1213 -815 -1147 -799
rect -1095 -765 -1029 -749
rect -1095 -799 -1079 -765
rect -1045 -799 -1029 -765
rect -1095 -815 -1029 -799
rect -977 -765 -911 -749
rect -977 -799 -961 -765
rect -927 -799 -911 -765
rect -977 -815 -911 -799
rect -859 -765 -793 -749
rect -859 -799 -843 -765
rect -809 -799 -793 -765
rect -859 -815 -793 -799
rect -741 -765 -675 -749
rect -741 -799 -725 -765
rect -691 -799 -675 -765
rect -741 -815 -675 -799
rect -623 -765 -557 -749
rect -623 -799 -607 -765
rect -573 -799 -557 -765
rect -623 -815 -557 -799
rect -505 -765 -439 -749
rect -505 -799 -489 -765
rect -455 -799 -439 -765
rect -505 -815 -439 -799
rect -387 -765 -321 -749
rect -387 -799 -371 -765
rect -337 -799 -321 -765
rect -387 -815 -321 -799
rect -269 -765 -203 -749
rect -269 -799 -253 -765
rect -219 -799 -203 -765
rect -269 -815 -203 -799
rect -151 -765 -85 -749
rect -151 -799 -135 -765
rect -101 -799 -85 -765
rect -151 -815 -85 -799
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect 85 -765 151 -749
rect 85 -799 101 -765
rect 135 -799 151 -765
rect 85 -815 151 -799
rect 203 -765 269 -749
rect 203 -799 219 -765
rect 253 -799 269 -765
rect 203 -815 269 -799
rect 321 -765 387 -749
rect 321 -799 337 -765
rect 371 -799 387 -765
rect 321 -815 387 -799
rect 439 -765 505 -749
rect 439 -799 455 -765
rect 489 -799 505 -765
rect 439 -815 505 -799
rect 557 -765 623 -749
rect 557 -799 573 -765
rect 607 -799 623 -765
rect 557 -815 623 -799
rect 675 -765 741 -749
rect 675 -799 691 -765
rect 725 -799 741 -765
rect 675 -815 741 -799
rect 793 -765 859 -749
rect 793 -799 809 -765
rect 843 -799 859 -765
rect 793 -815 859 -799
rect 911 -765 977 -749
rect 911 -799 927 -765
rect 961 -799 977 -765
rect 911 -815 977 -799
rect 1029 -765 1095 -749
rect 1029 -799 1045 -765
rect 1079 -799 1095 -765
rect 1029 -815 1095 -799
rect 1147 -765 1213 -749
rect 1147 -799 1163 -765
rect 1197 -799 1213 -765
rect 1147 -815 1213 -799
rect 1265 -765 1331 -749
rect 1265 -799 1281 -765
rect 1315 -799 1331 -765
rect 1265 -815 1331 -799
rect 1383 -765 1449 -749
rect 1383 -799 1399 -765
rect 1433 -799 1449 -765
rect 1383 -815 1449 -799
rect 1501 -765 1567 -749
rect 1501 -799 1517 -765
rect 1551 -799 1567 -765
rect 1501 -815 1567 -799
rect 1619 -765 1685 -749
rect 1619 -799 1635 -765
rect 1669 -799 1685 -765
rect 1619 -815 1685 -799
rect 1737 -765 1803 -749
rect 1737 -799 1753 -765
rect 1787 -799 1803 -765
rect 1737 -815 1803 -799
rect 1855 -765 1921 -749
rect 1855 -799 1871 -765
rect 1905 -799 1921 -765
rect 1855 -815 1921 -799
rect 1973 -765 2039 -749
rect 1973 -799 1989 -765
rect 2023 -799 2039 -765
rect 1973 -815 2039 -799
rect 2091 -765 2157 -749
rect 2091 -799 2107 -765
rect 2141 -799 2157 -765
rect 2091 -815 2157 -799
rect 2209 -765 2275 -749
rect 2209 -799 2225 -765
rect 2259 -799 2275 -765
rect 2209 -815 2275 -799
rect 2327 -765 2393 -749
rect 2327 -799 2343 -765
rect 2377 -799 2393 -765
rect 2327 -815 2393 -799
rect 2445 -765 2511 -749
rect 2445 -799 2461 -765
rect 2495 -799 2511 -765
rect 2445 -815 2511 -799
rect 2563 -765 2629 -749
rect 2563 -799 2579 -765
rect 2613 -799 2629 -765
rect 2563 -815 2629 -799
rect 2681 -765 2747 -749
rect 2681 -799 2697 -765
rect 2731 -799 2747 -765
rect 2681 -815 2747 -799
rect 2799 -765 2865 -749
rect 2799 -799 2815 -765
rect 2849 -799 2865 -765
rect 2799 -815 2865 -799
rect 2917 -765 2983 -749
rect 2917 -799 2933 -765
rect 2967 -799 2983 -765
rect 2917 -815 2983 -799
rect 3035 -765 3101 -749
rect 3035 -799 3051 -765
rect 3085 -799 3101 -765
rect 3035 -815 3101 -799
rect 3153 -765 3219 -749
rect 3153 -799 3169 -765
rect 3203 -799 3219 -765
rect 3153 -815 3219 -799
rect 3271 -765 3337 -749
rect 3271 -799 3287 -765
rect 3321 -799 3337 -765
rect 3271 -815 3337 -799
rect 3389 -765 3455 -749
rect 3389 -799 3405 -765
rect 3439 -799 3455 -765
rect 3389 -815 3455 -799
rect 3507 -765 3573 -749
rect 3507 -799 3523 -765
rect 3557 -799 3573 -765
rect 3507 -815 3573 -799
rect 3625 -765 3691 -749
rect 3625 -799 3641 -765
rect 3675 -799 3691 -765
rect 3625 -815 3691 -799
rect 3743 -765 3809 -749
rect 3743 -799 3759 -765
rect 3793 -799 3809 -765
rect 3743 -815 3809 -799
rect 3861 -765 3927 -749
rect 3861 -799 3877 -765
rect 3911 -799 3927 -765
rect 3861 -815 3927 -799
rect 3979 -765 4045 -749
rect 3979 -799 3995 -765
rect 4029 -799 4045 -765
rect 3979 -815 4045 -799
rect 4097 -765 4163 -749
rect 4097 -799 4113 -765
rect 4147 -799 4163 -765
rect 4097 -815 4163 -799
rect 4215 -765 4281 -749
rect 4215 -799 4231 -765
rect 4265 -799 4281 -765
rect 4215 -815 4281 -799
rect 4333 -765 4399 -749
rect 4333 -799 4349 -765
rect 4383 -799 4399 -765
rect 4333 -815 4399 -799
<< polycont >>
rect -4383 765 -4349 799
rect -4265 765 -4231 799
rect -4147 765 -4113 799
rect -4029 765 -3995 799
rect -3911 765 -3877 799
rect -3793 765 -3759 799
rect -3675 765 -3641 799
rect -3557 765 -3523 799
rect -3439 765 -3405 799
rect -3321 765 -3287 799
rect -3203 765 -3169 799
rect -3085 765 -3051 799
rect -2967 765 -2933 799
rect -2849 765 -2815 799
rect -2731 765 -2697 799
rect -2613 765 -2579 799
rect -2495 765 -2461 799
rect -2377 765 -2343 799
rect -2259 765 -2225 799
rect -2141 765 -2107 799
rect -2023 765 -1989 799
rect -1905 765 -1871 799
rect -1787 765 -1753 799
rect -1669 765 -1635 799
rect -1551 765 -1517 799
rect -1433 765 -1399 799
rect -1315 765 -1281 799
rect -1197 765 -1163 799
rect -1079 765 -1045 799
rect -961 765 -927 799
rect -843 765 -809 799
rect -725 765 -691 799
rect -607 765 -573 799
rect -489 765 -455 799
rect -371 765 -337 799
rect -253 765 -219 799
rect -135 765 -101 799
rect -17 765 17 799
rect 101 765 135 799
rect 219 765 253 799
rect 337 765 371 799
rect 455 765 489 799
rect 573 765 607 799
rect 691 765 725 799
rect 809 765 843 799
rect 927 765 961 799
rect 1045 765 1079 799
rect 1163 765 1197 799
rect 1281 765 1315 799
rect 1399 765 1433 799
rect 1517 765 1551 799
rect 1635 765 1669 799
rect 1753 765 1787 799
rect 1871 765 1905 799
rect 1989 765 2023 799
rect 2107 765 2141 799
rect 2225 765 2259 799
rect 2343 765 2377 799
rect 2461 765 2495 799
rect 2579 765 2613 799
rect 2697 765 2731 799
rect 2815 765 2849 799
rect 2933 765 2967 799
rect 3051 765 3085 799
rect 3169 765 3203 799
rect 3287 765 3321 799
rect 3405 765 3439 799
rect 3523 765 3557 799
rect 3641 765 3675 799
rect 3759 765 3793 799
rect 3877 765 3911 799
rect 3995 765 4029 799
rect 4113 765 4147 799
rect 4231 765 4265 799
rect 4349 765 4383 799
rect -4383 37 -4349 71
rect -4265 37 -4231 71
rect -4147 37 -4113 71
rect -4029 37 -3995 71
rect -3911 37 -3877 71
rect -3793 37 -3759 71
rect -3675 37 -3641 71
rect -3557 37 -3523 71
rect -3439 37 -3405 71
rect -3321 37 -3287 71
rect -3203 37 -3169 71
rect -3085 37 -3051 71
rect -2967 37 -2933 71
rect -2849 37 -2815 71
rect -2731 37 -2697 71
rect -2613 37 -2579 71
rect -2495 37 -2461 71
rect -2377 37 -2343 71
rect -2259 37 -2225 71
rect -2141 37 -2107 71
rect -2023 37 -1989 71
rect -1905 37 -1871 71
rect -1787 37 -1753 71
rect -1669 37 -1635 71
rect -1551 37 -1517 71
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect 1517 37 1551 71
rect 1635 37 1669 71
rect 1753 37 1787 71
rect 1871 37 1905 71
rect 1989 37 2023 71
rect 2107 37 2141 71
rect 2225 37 2259 71
rect 2343 37 2377 71
rect 2461 37 2495 71
rect 2579 37 2613 71
rect 2697 37 2731 71
rect 2815 37 2849 71
rect 2933 37 2967 71
rect 3051 37 3085 71
rect 3169 37 3203 71
rect 3287 37 3321 71
rect 3405 37 3439 71
rect 3523 37 3557 71
rect 3641 37 3675 71
rect 3759 37 3793 71
rect 3877 37 3911 71
rect 3995 37 4029 71
rect 4113 37 4147 71
rect 4231 37 4265 71
rect 4349 37 4383 71
rect -4383 -71 -4349 -37
rect -4265 -71 -4231 -37
rect -4147 -71 -4113 -37
rect -4029 -71 -3995 -37
rect -3911 -71 -3877 -37
rect -3793 -71 -3759 -37
rect -3675 -71 -3641 -37
rect -3557 -71 -3523 -37
rect -3439 -71 -3405 -37
rect -3321 -71 -3287 -37
rect -3203 -71 -3169 -37
rect -3085 -71 -3051 -37
rect -2967 -71 -2933 -37
rect -2849 -71 -2815 -37
rect -2731 -71 -2697 -37
rect -2613 -71 -2579 -37
rect -2495 -71 -2461 -37
rect -2377 -71 -2343 -37
rect -2259 -71 -2225 -37
rect -2141 -71 -2107 -37
rect -2023 -71 -1989 -37
rect -1905 -71 -1871 -37
rect -1787 -71 -1753 -37
rect -1669 -71 -1635 -37
rect -1551 -71 -1517 -37
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
rect 1517 -71 1551 -37
rect 1635 -71 1669 -37
rect 1753 -71 1787 -37
rect 1871 -71 1905 -37
rect 1989 -71 2023 -37
rect 2107 -71 2141 -37
rect 2225 -71 2259 -37
rect 2343 -71 2377 -37
rect 2461 -71 2495 -37
rect 2579 -71 2613 -37
rect 2697 -71 2731 -37
rect 2815 -71 2849 -37
rect 2933 -71 2967 -37
rect 3051 -71 3085 -37
rect 3169 -71 3203 -37
rect 3287 -71 3321 -37
rect 3405 -71 3439 -37
rect 3523 -71 3557 -37
rect 3641 -71 3675 -37
rect 3759 -71 3793 -37
rect 3877 -71 3911 -37
rect 3995 -71 4029 -37
rect 4113 -71 4147 -37
rect 4231 -71 4265 -37
rect 4349 -71 4383 -37
rect -4383 -799 -4349 -765
rect -4265 -799 -4231 -765
rect -4147 -799 -4113 -765
rect -4029 -799 -3995 -765
rect -3911 -799 -3877 -765
rect -3793 -799 -3759 -765
rect -3675 -799 -3641 -765
rect -3557 -799 -3523 -765
rect -3439 -799 -3405 -765
rect -3321 -799 -3287 -765
rect -3203 -799 -3169 -765
rect -3085 -799 -3051 -765
rect -2967 -799 -2933 -765
rect -2849 -799 -2815 -765
rect -2731 -799 -2697 -765
rect -2613 -799 -2579 -765
rect -2495 -799 -2461 -765
rect -2377 -799 -2343 -765
rect -2259 -799 -2225 -765
rect -2141 -799 -2107 -765
rect -2023 -799 -1989 -765
rect -1905 -799 -1871 -765
rect -1787 -799 -1753 -765
rect -1669 -799 -1635 -765
rect -1551 -799 -1517 -765
rect -1433 -799 -1399 -765
rect -1315 -799 -1281 -765
rect -1197 -799 -1163 -765
rect -1079 -799 -1045 -765
rect -961 -799 -927 -765
rect -843 -799 -809 -765
rect -725 -799 -691 -765
rect -607 -799 -573 -765
rect -489 -799 -455 -765
rect -371 -799 -337 -765
rect -253 -799 -219 -765
rect -135 -799 -101 -765
rect -17 -799 17 -765
rect 101 -799 135 -765
rect 219 -799 253 -765
rect 337 -799 371 -765
rect 455 -799 489 -765
rect 573 -799 607 -765
rect 691 -799 725 -765
rect 809 -799 843 -765
rect 927 -799 961 -765
rect 1045 -799 1079 -765
rect 1163 -799 1197 -765
rect 1281 -799 1315 -765
rect 1399 -799 1433 -765
rect 1517 -799 1551 -765
rect 1635 -799 1669 -765
rect 1753 -799 1787 -765
rect 1871 -799 1905 -765
rect 1989 -799 2023 -765
rect 2107 -799 2141 -765
rect 2225 -799 2259 -765
rect 2343 -799 2377 -765
rect 2461 -799 2495 -765
rect 2579 -799 2613 -765
rect 2697 -799 2731 -765
rect 2815 -799 2849 -765
rect 2933 -799 2967 -765
rect 3051 -799 3085 -765
rect 3169 -799 3203 -765
rect 3287 -799 3321 -765
rect 3405 -799 3439 -765
rect 3523 -799 3557 -765
rect 3641 -799 3675 -765
rect 3759 -799 3793 -765
rect 3877 -799 3911 -765
rect 3995 -799 4029 -765
rect 4113 -799 4147 -765
rect 4231 -799 4265 -765
rect 4349 -799 4383 -765
<< locali >>
rect -4556 867 -4460 901
rect 4460 867 4556 901
rect -4556 805 -4522 867
rect 4522 805 4556 867
rect -4399 765 -4383 799
rect -4349 765 -4333 799
rect -4281 765 -4265 799
rect -4231 765 -4215 799
rect -4163 765 -4147 799
rect -4113 765 -4097 799
rect -4045 765 -4029 799
rect -3995 765 -3979 799
rect -3927 765 -3911 799
rect -3877 765 -3861 799
rect -3809 765 -3793 799
rect -3759 765 -3743 799
rect -3691 765 -3675 799
rect -3641 765 -3625 799
rect -3573 765 -3557 799
rect -3523 765 -3507 799
rect -3455 765 -3439 799
rect -3405 765 -3389 799
rect -3337 765 -3321 799
rect -3287 765 -3271 799
rect -3219 765 -3203 799
rect -3169 765 -3153 799
rect -3101 765 -3085 799
rect -3051 765 -3035 799
rect -2983 765 -2967 799
rect -2933 765 -2917 799
rect -2865 765 -2849 799
rect -2815 765 -2799 799
rect -2747 765 -2731 799
rect -2697 765 -2681 799
rect -2629 765 -2613 799
rect -2579 765 -2563 799
rect -2511 765 -2495 799
rect -2461 765 -2445 799
rect -2393 765 -2377 799
rect -2343 765 -2327 799
rect -2275 765 -2259 799
rect -2225 765 -2209 799
rect -2157 765 -2141 799
rect -2107 765 -2091 799
rect -2039 765 -2023 799
rect -1989 765 -1973 799
rect -1921 765 -1905 799
rect -1871 765 -1855 799
rect -1803 765 -1787 799
rect -1753 765 -1737 799
rect -1685 765 -1669 799
rect -1635 765 -1619 799
rect -1567 765 -1551 799
rect -1517 765 -1501 799
rect -1449 765 -1433 799
rect -1399 765 -1383 799
rect -1331 765 -1315 799
rect -1281 765 -1265 799
rect -1213 765 -1197 799
rect -1163 765 -1147 799
rect -1095 765 -1079 799
rect -1045 765 -1029 799
rect -977 765 -961 799
rect -927 765 -911 799
rect -859 765 -843 799
rect -809 765 -793 799
rect -741 765 -725 799
rect -691 765 -675 799
rect -623 765 -607 799
rect -573 765 -557 799
rect -505 765 -489 799
rect -455 765 -439 799
rect -387 765 -371 799
rect -337 765 -321 799
rect -269 765 -253 799
rect -219 765 -203 799
rect -151 765 -135 799
rect -101 765 -85 799
rect -33 765 -17 799
rect 17 765 33 799
rect 85 765 101 799
rect 135 765 151 799
rect 203 765 219 799
rect 253 765 269 799
rect 321 765 337 799
rect 371 765 387 799
rect 439 765 455 799
rect 489 765 505 799
rect 557 765 573 799
rect 607 765 623 799
rect 675 765 691 799
rect 725 765 741 799
rect 793 765 809 799
rect 843 765 859 799
rect 911 765 927 799
rect 961 765 977 799
rect 1029 765 1045 799
rect 1079 765 1095 799
rect 1147 765 1163 799
rect 1197 765 1213 799
rect 1265 765 1281 799
rect 1315 765 1331 799
rect 1383 765 1399 799
rect 1433 765 1449 799
rect 1501 765 1517 799
rect 1551 765 1567 799
rect 1619 765 1635 799
rect 1669 765 1685 799
rect 1737 765 1753 799
rect 1787 765 1803 799
rect 1855 765 1871 799
rect 1905 765 1921 799
rect 1973 765 1989 799
rect 2023 765 2039 799
rect 2091 765 2107 799
rect 2141 765 2157 799
rect 2209 765 2225 799
rect 2259 765 2275 799
rect 2327 765 2343 799
rect 2377 765 2393 799
rect 2445 765 2461 799
rect 2495 765 2511 799
rect 2563 765 2579 799
rect 2613 765 2629 799
rect 2681 765 2697 799
rect 2731 765 2747 799
rect 2799 765 2815 799
rect 2849 765 2865 799
rect 2917 765 2933 799
rect 2967 765 2983 799
rect 3035 765 3051 799
rect 3085 765 3101 799
rect 3153 765 3169 799
rect 3203 765 3219 799
rect 3271 765 3287 799
rect 3321 765 3337 799
rect 3389 765 3405 799
rect 3439 765 3455 799
rect 3507 765 3523 799
rect 3557 765 3573 799
rect 3625 765 3641 799
rect 3675 765 3691 799
rect 3743 765 3759 799
rect 3793 765 3809 799
rect 3861 765 3877 799
rect 3911 765 3927 799
rect 3979 765 3995 799
rect 4029 765 4045 799
rect 4097 765 4113 799
rect 4147 765 4163 799
rect 4215 765 4231 799
rect 4265 765 4281 799
rect 4333 765 4349 799
rect 4383 765 4399 799
rect -4442 706 -4408 722
rect -4442 114 -4408 130
rect -4324 706 -4290 722
rect -4324 114 -4290 130
rect -4206 706 -4172 722
rect -4206 114 -4172 130
rect -4088 706 -4054 722
rect -4088 114 -4054 130
rect -3970 706 -3936 722
rect -3970 114 -3936 130
rect -3852 706 -3818 722
rect -3852 114 -3818 130
rect -3734 706 -3700 722
rect -3734 114 -3700 130
rect -3616 706 -3582 722
rect -3616 114 -3582 130
rect -3498 706 -3464 722
rect -3498 114 -3464 130
rect -3380 706 -3346 722
rect -3380 114 -3346 130
rect -3262 706 -3228 722
rect -3262 114 -3228 130
rect -3144 706 -3110 722
rect -3144 114 -3110 130
rect -3026 706 -2992 722
rect -3026 114 -2992 130
rect -2908 706 -2874 722
rect -2908 114 -2874 130
rect -2790 706 -2756 722
rect -2790 114 -2756 130
rect -2672 706 -2638 722
rect -2672 114 -2638 130
rect -2554 706 -2520 722
rect -2554 114 -2520 130
rect -2436 706 -2402 722
rect -2436 114 -2402 130
rect -2318 706 -2284 722
rect -2318 114 -2284 130
rect -2200 706 -2166 722
rect -2200 114 -2166 130
rect -2082 706 -2048 722
rect -2082 114 -2048 130
rect -1964 706 -1930 722
rect -1964 114 -1930 130
rect -1846 706 -1812 722
rect -1846 114 -1812 130
rect -1728 706 -1694 722
rect -1728 114 -1694 130
rect -1610 706 -1576 722
rect -1610 114 -1576 130
rect -1492 706 -1458 722
rect -1492 114 -1458 130
rect -1374 706 -1340 722
rect -1374 114 -1340 130
rect -1256 706 -1222 722
rect -1256 114 -1222 130
rect -1138 706 -1104 722
rect -1138 114 -1104 130
rect -1020 706 -986 722
rect -1020 114 -986 130
rect -902 706 -868 722
rect -902 114 -868 130
rect -784 706 -750 722
rect -784 114 -750 130
rect -666 706 -632 722
rect -666 114 -632 130
rect -548 706 -514 722
rect -548 114 -514 130
rect -430 706 -396 722
rect -430 114 -396 130
rect -312 706 -278 722
rect -312 114 -278 130
rect -194 706 -160 722
rect -194 114 -160 130
rect -76 706 -42 722
rect -76 114 -42 130
rect 42 706 76 722
rect 42 114 76 130
rect 160 706 194 722
rect 160 114 194 130
rect 278 706 312 722
rect 278 114 312 130
rect 396 706 430 722
rect 396 114 430 130
rect 514 706 548 722
rect 514 114 548 130
rect 632 706 666 722
rect 632 114 666 130
rect 750 706 784 722
rect 750 114 784 130
rect 868 706 902 722
rect 868 114 902 130
rect 986 706 1020 722
rect 986 114 1020 130
rect 1104 706 1138 722
rect 1104 114 1138 130
rect 1222 706 1256 722
rect 1222 114 1256 130
rect 1340 706 1374 722
rect 1340 114 1374 130
rect 1458 706 1492 722
rect 1458 114 1492 130
rect 1576 706 1610 722
rect 1576 114 1610 130
rect 1694 706 1728 722
rect 1694 114 1728 130
rect 1812 706 1846 722
rect 1812 114 1846 130
rect 1930 706 1964 722
rect 1930 114 1964 130
rect 2048 706 2082 722
rect 2048 114 2082 130
rect 2166 706 2200 722
rect 2166 114 2200 130
rect 2284 706 2318 722
rect 2284 114 2318 130
rect 2402 706 2436 722
rect 2402 114 2436 130
rect 2520 706 2554 722
rect 2520 114 2554 130
rect 2638 706 2672 722
rect 2638 114 2672 130
rect 2756 706 2790 722
rect 2756 114 2790 130
rect 2874 706 2908 722
rect 2874 114 2908 130
rect 2992 706 3026 722
rect 2992 114 3026 130
rect 3110 706 3144 722
rect 3110 114 3144 130
rect 3228 706 3262 722
rect 3228 114 3262 130
rect 3346 706 3380 722
rect 3346 114 3380 130
rect 3464 706 3498 722
rect 3464 114 3498 130
rect 3582 706 3616 722
rect 3582 114 3616 130
rect 3700 706 3734 722
rect 3700 114 3734 130
rect 3818 706 3852 722
rect 3818 114 3852 130
rect 3936 706 3970 722
rect 3936 114 3970 130
rect 4054 706 4088 722
rect 4054 114 4088 130
rect 4172 706 4206 722
rect 4172 114 4206 130
rect 4290 706 4324 722
rect 4290 114 4324 130
rect 4408 706 4442 722
rect 4408 114 4442 130
rect -4399 37 -4383 71
rect -4349 37 -4333 71
rect -4281 37 -4265 71
rect -4231 37 -4215 71
rect -4163 37 -4147 71
rect -4113 37 -4097 71
rect -4045 37 -4029 71
rect -3995 37 -3979 71
rect -3927 37 -3911 71
rect -3877 37 -3861 71
rect -3809 37 -3793 71
rect -3759 37 -3743 71
rect -3691 37 -3675 71
rect -3641 37 -3625 71
rect -3573 37 -3557 71
rect -3523 37 -3507 71
rect -3455 37 -3439 71
rect -3405 37 -3389 71
rect -3337 37 -3321 71
rect -3287 37 -3271 71
rect -3219 37 -3203 71
rect -3169 37 -3153 71
rect -3101 37 -3085 71
rect -3051 37 -3035 71
rect -2983 37 -2967 71
rect -2933 37 -2917 71
rect -2865 37 -2849 71
rect -2815 37 -2799 71
rect -2747 37 -2731 71
rect -2697 37 -2681 71
rect -2629 37 -2613 71
rect -2579 37 -2563 71
rect -2511 37 -2495 71
rect -2461 37 -2445 71
rect -2393 37 -2377 71
rect -2343 37 -2327 71
rect -2275 37 -2259 71
rect -2225 37 -2209 71
rect -2157 37 -2141 71
rect -2107 37 -2091 71
rect -2039 37 -2023 71
rect -1989 37 -1973 71
rect -1921 37 -1905 71
rect -1871 37 -1855 71
rect -1803 37 -1787 71
rect -1753 37 -1737 71
rect -1685 37 -1669 71
rect -1635 37 -1619 71
rect -1567 37 -1551 71
rect -1517 37 -1501 71
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -977 37 -961 71
rect -927 37 -911 71
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect 911 37 927 71
rect 961 37 977 71
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1501 37 1517 71
rect 1551 37 1567 71
rect 1619 37 1635 71
rect 1669 37 1685 71
rect 1737 37 1753 71
rect 1787 37 1803 71
rect 1855 37 1871 71
rect 1905 37 1921 71
rect 1973 37 1989 71
rect 2023 37 2039 71
rect 2091 37 2107 71
rect 2141 37 2157 71
rect 2209 37 2225 71
rect 2259 37 2275 71
rect 2327 37 2343 71
rect 2377 37 2393 71
rect 2445 37 2461 71
rect 2495 37 2511 71
rect 2563 37 2579 71
rect 2613 37 2629 71
rect 2681 37 2697 71
rect 2731 37 2747 71
rect 2799 37 2815 71
rect 2849 37 2865 71
rect 2917 37 2933 71
rect 2967 37 2983 71
rect 3035 37 3051 71
rect 3085 37 3101 71
rect 3153 37 3169 71
rect 3203 37 3219 71
rect 3271 37 3287 71
rect 3321 37 3337 71
rect 3389 37 3405 71
rect 3439 37 3455 71
rect 3507 37 3523 71
rect 3557 37 3573 71
rect 3625 37 3641 71
rect 3675 37 3691 71
rect 3743 37 3759 71
rect 3793 37 3809 71
rect 3861 37 3877 71
rect 3911 37 3927 71
rect 3979 37 3995 71
rect 4029 37 4045 71
rect 4097 37 4113 71
rect 4147 37 4163 71
rect 4215 37 4231 71
rect 4265 37 4281 71
rect 4333 37 4349 71
rect 4383 37 4399 71
rect -4399 -71 -4383 -37
rect -4349 -71 -4333 -37
rect -4281 -71 -4265 -37
rect -4231 -71 -4215 -37
rect -4163 -71 -4147 -37
rect -4113 -71 -4097 -37
rect -4045 -71 -4029 -37
rect -3995 -71 -3979 -37
rect -3927 -71 -3911 -37
rect -3877 -71 -3861 -37
rect -3809 -71 -3793 -37
rect -3759 -71 -3743 -37
rect -3691 -71 -3675 -37
rect -3641 -71 -3625 -37
rect -3573 -71 -3557 -37
rect -3523 -71 -3507 -37
rect -3455 -71 -3439 -37
rect -3405 -71 -3389 -37
rect -3337 -71 -3321 -37
rect -3287 -71 -3271 -37
rect -3219 -71 -3203 -37
rect -3169 -71 -3153 -37
rect -3101 -71 -3085 -37
rect -3051 -71 -3035 -37
rect -2983 -71 -2967 -37
rect -2933 -71 -2917 -37
rect -2865 -71 -2849 -37
rect -2815 -71 -2799 -37
rect -2747 -71 -2731 -37
rect -2697 -71 -2681 -37
rect -2629 -71 -2613 -37
rect -2579 -71 -2563 -37
rect -2511 -71 -2495 -37
rect -2461 -71 -2445 -37
rect -2393 -71 -2377 -37
rect -2343 -71 -2327 -37
rect -2275 -71 -2259 -37
rect -2225 -71 -2209 -37
rect -2157 -71 -2141 -37
rect -2107 -71 -2091 -37
rect -2039 -71 -2023 -37
rect -1989 -71 -1973 -37
rect -1921 -71 -1905 -37
rect -1871 -71 -1855 -37
rect -1803 -71 -1787 -37
rect -1753 -71 -1737 -37
rect -1685 -71 -1669 -37
rect -1635 -71 -1619 -37
rect -1567 -71 -1551 -37
rect -1517 -71 -1501 -37
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect 1501 -71 1517 -37
rect 1551 -71 1567 -37
rect 1619 -71 1635 -37
rect 1669 -71 1685 -37
rect 1737 -71 1753 -37
rect 1787 -71 1803 -37
rect 1855 -71 1871 -37
rect 1905 -71 1921 -37
rect 1973 -71 1989 -37
rect 2023 -71 2039 -37
rect 2091 -71 2107 -37
rect 2141 -71 2157 -37
rect 2209 -71 2225 -37
rect 2259 -71 2275 -37
rect 2327 -71 2343 -37
rect 2377 -71 2393 -37
rect 2445 -71 2461 -37
rect 2495 -71 2511 -37
rect 2563 -71 2579 -37
rect 2613 -71 2629 -37
rect 2681 -71 2697 -37
rect 2731 -71 2747 -37
rect 2799 -71 2815 -37
rect 2849 -71 2865 -37
rect 2917 -71 2933 -37
rect 2967 -71 2983 -37
rect 3035 -71 3051 -37
rect 3085 -71 3101 -37
rect 3153 -71 3169 -37
rect 3203 -71 3219 -37
rect 3271 -71 3287 -37
rect 3321 -71 3337 -37
rect 3389 -71 3405 -37
rect 3439 -71 3455 -37
rect 3507 -71 3523 -37
rect 3557 -71 3573 -37
rect 3625 -71 3641 -37
rect 3675 -71 3691 -37
rect 3743 -71 3759 -37
rect 3793 -71 3809 -37
rect 3861 -71 3877 -37
rect 3911 -71 3927 -37
rect 3979 -71 3995 -37
rect 4029 -71 4045 -37
rect 4097 -71 4113 -37
rect 4147 -71 4163 -37
rect 4215 -71 4231 -37
rect 4265 -71 4281 -37
rect 4333 -71 4349 -37
rect 4383 -71 4399 -37
rect -4442 -130 -4408 -114
rect -4442 -722 -4408 -706
rect -4324 -130 -4290 -114
rect -4324 -722 -4290 -706
rect -4206 -130 -4172 -114
rect -4206 -722 -4172 -706
rect -4088 -130 -4054 -114
rect -4088 -722 -4054 -706
rect -3970 -130 -3936 -114
rect -3970 -722 -3936 -706
rect -3852 -130 -3818 -114
rect -3852 -722 -3818 -706
rect -3734 -130 -3700 -114
rect -3734 -722 -3700 -706
rect -3616 -130 -3582 -114
rect -3616 -722 -3582 -706
rect -3498 -130 -3464 -114
rect -3498 -722 -3464 -706
rect -3380 -130 -3346 -114
rect -3380 -722 -3346 -706
rect -3262 -130 -3228 -114
rect -3262 -722 -3228 -706
rect -3144 -130 -3110 -114
rect -3144 -722 -3110 -706
rect -3026 -130 -2992 -114
rect -3026 -722 -2992 -706
rect -2908 -130 -2874 -114
rect -2908 -722 -2874 -706
rect -2790 -130 -2756 -114
rect -2790 -722 -2756 -706
rect -2672 -130 -2638 -114
rect -2672 -722 -2638 -706
rect -2554 -130 -2520 -114
rect -2554 -722 -2520 -706
rect -2436 -130 -2402 -114
rect -2436 -722 -2402 -706
rect -2318 -130 -2284 -114
rect -2318 -722 -2284 -706
rect -2200 -130 -2166 -114
rect -2200 -722 -2166 -706
rect -2082 -130 -2048 -114
rect -2082 -722 -2048 -706
rect -1964 -130 -1930 -114
rect -1964 -722 -1930 -706
rect -1846 -130 -1812 -114
rect -1846 -722 -1812 -706
rect -1728 -130 -1694 -114
rect -1728 -722 -1694 -706
rect -1610 -130 -1576 -114
rect -1610 -722 -1576 -706
rect -1492 -130 -1458 -114
rect -1492 -722 -1458 -706
rect -1374 -130 -1340 -114
rect -1374 -722 -1340 -706
rect -1256 -130 -1222 -114
rect -1256 -722 -1222 -706
rect -1138 -130 -1104 -114
rect -1138 -722 -1104 -706
rect -1020 -130 -986 -114
rect -1020 -722 -986 -706
rect -902 -130 -868 -114
rect -902 -722 -868 -706
rect -784 -130 -750 -114
rect -784 -722 -750 -706
rect -666 -130 -632 -114
rect -666 -722 -632 -706
rect -548 -130 -514 -114
rect -548 -722 -514 -706
rect -430 -130 -396 -114
rect -430 -722 -396 -706
rect -312 -130 -278 -114
rect -312 -722 -278 -706
rect -194 -130 -160 -114
rect -194 -722 -160 -706
rect -76 -130 -42 -114
rect -76 -722 -42 -706
rect 42 -130 76 -114
rect 42 -722 76 -706
rect 160 -130 194 -114
rect 160 -722 194 -706
rect 278 -130 312 -114
rect 278 -722 312 -706
rect 396 -130 430 -114
rect 396 -722 430 -706
rect 514 -130 548 -114
rect 514 -722 548 -706
rect 632 -130 666 -114
rect 632 -722 666 -706
rect 750 -130 784 -114
rect 750 -722 784 -706
rect 868 -130 902 -114
rect 868 -722 902 -706
rect 986 -130 1020 -114
rect 986 -722 1020 -706
rect 1104 -130 1138 -114
rect 1104 -722 1138 -706
rect 1222 -130 1256 -114
rect 1222 -722 1256 -706
rect 1340 -130 1374 -114
rect 1340 -722 1374 -706
rect 1458 -130 1492 -114
rect 1458 -722 1492 -706
rect 1576 -130 1610 -114
rect 1576 -722 1610 -706
rect 1694 -130 1728 -114
rect 1694 -722 1728 -706
rect 1812 -130 1846 -114
rect 1812 -722 1846 -706
rect 1930 -130 1964 -114
rect 1930 -722 1964 -706
rect 2048 -130 2082 -114
rect 2048 -722 2082 -706
rect 2166 -130 2200 -114
rect 2166 -722 2200 -706
rect 2284 -130 2318 -114
rect 2284 -722 2318 -706
rect 2402 -130 2436 -114
rect 2402 -722 2436 -706
rect 2520 -130 2554 -114
rect 2520 -722 2554 -706
rect 2638 -130 2672 -114
rect 2638 -722 2672 -706
rect 2756 -130 2790 -114
rect 2756 -722 2790 -706
rect 2874 -130 2908 -114
rect 2874 -722 2908 -706
rect 2992 -130 3026 -114
rect 2992 -722 3026 -706
rect 3110 -130 3144 -114
rect 3110 -722 3144 -706
rect 3228 -130 3262 -114
rect 3228 -722 3262 -706
rect 3346 -130 3380 -114
rect 3346 -722 3380 -706
rect 3464 -130 3498 -114
rect 3464 -722 3498 -706
rect 3582 -130 3616 -114
rect 3582 -722 3616 -706
rect 3700 -130 3734 -114
rect 3700 -722 3734 -706
rect 3818 -130 3852 -114
rect 3818 -722 3852 -706
rect 3936 -130 3970 -114
rect 3936 -722 3970 -706
rect 4054 -130 4088 -114
rect 4054 -722 4088 -706
rect 4172 -130 4206 -114
rect 4172 -722 4206 -706
rect 4290 -130 4324 -114
rect 4290 -722 4324 -706
rect 4408 -130 4442 -114
rect 4408 -722 4442 -706
rect -4399 -799 -4383 -765
rect -4349 -799 -4333 -765
rect -4281 -799 -4265 -765
rect -4231 -799 -4215 -765
rect -4163 -799 -4147 -765
rect -4113 -799 -4097 -765
rect -4045 -799 -4029 -765
rect -3995 -799 -3979 -765
rect -3927 -799 -3911 -765
rect -3877 -799 -3861 -765
rect -3809 -799 -3793 -765
rect -3759 -799 -3743 -765
rect -3691 -799 -3675 -765
rect -3641 -799 -3625 -765
rect -3573 -799 -3557 -765
rect -3523 -799 -3507 -765
rect -3455 -799 -3439 -765
rect -3405 -799 -3389 -765
rect -3337 -799 -3321 -765
rect -3287 -799 -3271 -765
rect -3219 -799 -3203 -765
rect -3169 -799 -3153 -765
rect -3101 -799 -3085 -765
rect -3051 -799 -3035 -765
rect -2983 -799 -2967 -765
rect -2933 -799 -2917 -765
rect -2865 -799 -2849 -765
rect -2815 -799 -2799 -765
rect -2747 -799 -2731 -765
rect -2697 -799 -2681 -765
rect -2629 -799 -2613 -765
rect -2579 -799 -2563 -765
rect -2511 -799 -2495 -765
rect -2461 -799 -2445 -765
rect -2393 -799 -2377 -765
rect -2343 -799 -2327 -765
rect -2275 -799 -2259 -765
rect -2225 -799 -2209 -765
rect -2157 -799 -2141 -765
rect -2107 -799 -2091 -765
rect -2039 -799 -2023 -765
rect -1989 -799 -1973 -765
rect -1921 -799 -1905 -765
rect -1871 -799 -1855 -765
rect -1803 -799 -1787 -765
rect -1753 -799 -1737 -765
rect -1685 -799 -1669 -765
rect -1635 -799 -1619 -765
rect -1567 -799 -1551 -765
rect -1517 -799 -1501 -765
rect -1449 -799 -1433 -765
rect -1399 -799 -1383 -765
rect -1331 -799 -1315 -765
rect -1281 -799 -1265 -765
rect -1213 -799 -1197 -765
rect -1163 -799 -1147 -765
rect -1095 -799 -1079 -765
rect -1045 -799 -1029 -765
rect -977 -799 -961 -765
rect -927 -799 -911 -765
rect -859 -799 -843 -765
rect -809 -799 -793 -765
rect -741 -799 -725 -765
rect -691 -799 -675 -765
rect -623 -799 -607 -765
rect -573 -799 -557 -765
rect -505 -799 -489 -765
rect -455 -799 -439 -765
rect -387 -799 -371 -765
rect -337 -799 -321 -765
rect -269 -799 -253 -765
rect -219 -799 -203 -765
rect -151 -799 -135 -765
rect -101 -799 -85 -765
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect 85 -799 101 -765
rect 135 -799 151 -765
rect 203 -799 219 -765
rect 253 -799 269 -765
rect 321 -799 337 -765
rect 371 -799 387 -765
rect 439 -799 455 -765
rect 489 -799 505 -765
rect 557 -799 573 -765
rect 607 -799 623 -765
rect 675 -799 691 -765
rect 725 -799 741 -765
rect 793 -799 809 -765
rect 843 -799 859 -765
rect 911 -799 927 -765
rect 961 -799 977 -765
rect 1029 -799 1045 -765
rect 1079 -799 1095 -765
rect 1147 -799 1163 -765
rect 1197 -799 1213 -765
rect 1265 -799 1281 -765
rect 1315 -799 1331 -765
rect 1383 -799 1399 -765
rect 1433 -799 1449 -765
rect 1501 -799 1517 -765
rect 1551 -799 1567 -765
rect 1619 -799 1635 -765
rect 1669 -799 1685 -765
rect 1737 -799 1753 -765
rect 1787 -799 1803 -765
rect 1855 -799 1871 -765
rect 1905 -799 1921 -765
rect 1973 -799 1989 -765
rect 2023 -799 2039 -765
rect 2091 -799 2107 -765
rect 2141 -799 2157 -765
rect 2209 -799 2225 -765
rect 2259 -799 2275 -765
rect 2327 -799 2343 -765
rect 2377 -799 2393 -765
rect 2445 -799 2461 -765
rect 2495 -799 2511 -765
rect 2563 -799 2579 -765
rect 2613 -799 2629 -765
rect 2681 -799 2697 -765
rect 2731 -799 2747 -765
rect 2799 -799 2815 -765
rect 2849 -799 2865 -765
rect 2917 -799 2933 -765
rect 2967 -799 2983 -765
rect 3035 -799 3051 -765
rect 3085 -799 3101 -765
rect 3153 -799 3169 -765
rect 3203 -799 3219 -765
rect 3271 -799 3287 -765
rect 3321 -799 3337 -765
rect 3389 -799 3405 -765
rect 3439 -799 3455 -765
rect 3507 -799 3523 -765
rect 3557 -799 3573 -765
rect 3625 -799 3641 -765
rect 3675 -799 3691 -765
rect 3743 -799 3759 -765
rect 3793 -799 3809 -765
rect 3861 -799 3877 -765
rect 3911 -799 3927 -765
rect 3979 -799 3995 -765
rect 4029 -799 4045 -765
rect 4097 -799 4113 -765
rect 4147 -799 4163 -765
rect 4215 -799 4231 -765
rect 4265 -799 4281 -765
rect 4333 -799 4349 -765
rect 4383 -799 4399 -765
rect -4556 -867 -4522 -805
rect 4522 -867 4556 -805
rect -4556 -901 -4460 -867
rect 4460 -901 4556 -867
<< viali >>
rect -4383 765 -4349 799
rect -4265 765 -4231 799
rect -4147 765 -4113 799
rect -4029 765 -3995 799
rect -3911 765 -3877 799
rect -3793 765 -3759 799
rect -3675 765 -3641 799
rect -3557 765 -3523 799
rect -3439 765 -3405 799
rect -3321 765 -3287 799
rect -3203 765 -3169 799
rect -3085 765 -3051 799
rect -2967 765 -2933 799
rect -2849 765 -2815 799
rect -2731 765 -2697 799
rect -2613 765 -2579 799
rect -2495 765 -2461 799
rect -2377 765 -2343 799
rect -2259 765 -2225 799
rect -2141 765 -2107 799
rect -2023 765 -1989 799
rect -1905 765 -1871 799
rect -1787 765 -1753 799
rect -1669 765 -1635 799
rect -1551 765 -1517 799
rect -1433 765 -1399 799
rect -1315 765 -1281 799
rect -1197 765 -1163 799
rect -1079 765 -1045 799
rect -961 765 -927 799
rect -843 765 -809 799
rect -725 765 -691 799
rect -607 765 -573 799
rect -489 765 -455 799
rect -371 765 -337 799
rect -253 765 -219 799
rect -135 765 -101 799
rect -17 765 17 799
rect 101 765 135 799
rect 219 765 253 799
rect 337 765 371 799
rect 455 765 489 799
rect 573 765 607 799
rect 691 765 725 799
rect 809 765 843 799
rect 927 765 961 799
rect 1045 765 1079 799
rect 1163 765 1197 799
rect 1281 765 1315 799
rect 1399 765 1433 799
rect 1517 765 1551 799
rect 1635 765 1669 799
rect 1753 765 1787 799
rect 1871 765 1905 799
rect 1989 765 2023 799
rect 2107 765 2141 799
rect 2225 765 2259 799
rect 2343 765 2377 799
rect 2461 765 2495 799
rect 2579 765 2613 799
rect 2697 765 2731 799
rect 2815 765 2849 799
rect 2933 765 2967 799
rect 3051 765 3085 799
rect 3169 765 3203 799
rect 3287 765 3321 799
rect 3405 765 3439 799
rect 3523 765 3557 799
rect 3641 765 3675 799
rect 3759 765 3793 799
rect 3877 765 3911 799
rect 3995 765 4029 799
rect 4113 765 4147 799
rect 4231 765 4265 799
rect 4349 765 4383 799
rect -4442 130 -4408 706
rect -4324 130 -4290 706
rect -4206 130 -4172 706
rect -4088 130 -4054 706
rect -3970 130 -3936 706
rect -3852 130 -3818 706
rect -3734 130 -3700 706
rect -3616 130 -3582 706
rect -3498 130 -3464 706
rect -3380 130 -3346 706
rect -3262 130 -3228 706
rect -3144 130 -3110 706
rect -3026 130 -2992 706
rect -2908 130 -2874 706
rect -2790 130 -2756 706
rect -2672 130 -2638 706
rect -2554 130 -2520 706
rect -2436 130 -2402 706
rect -2318 130 -2284 706
rect -2200 130 -2166 706
rect -2082 130 -2048 706
rect -1964 130 -1930 706
rect -1846 130 -1812 706
rect -1728 130 -1694 706
rect -1610 130 -1576 706
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect 1576 130 1610 706
rect 1694 130 1728 706
rect 1812 130 1846 706
rect 1930 130 1964 706
rect 2048 130 2082 706
rect 2166 130 2200 706
rect 2284 130 2318 706
rect 2402 130 2436 706
rect 2520 130 2554 706
rect 2638 130 2672 706
rect 2756 130 2790 706
rect 2874 130 2908 706
rect 2992 130 3026 706
rect 3110 130 3144 706
rect 3228 130 3262 706
rect 3346 130 3380 706
rect 3464 130 3498 706
rect 3582 130 3616 706
rect 3700 130 3734 706
rect 3818 130 3852 706
rect 3936 130 3970 706
rect 4054 130 4088 706
rect 4172 130 4206 706
rect 4290 130 4324 706
rect 4408 130 4442 706
rect -4383 37 -4349 71
rect -4265 37 -4231 71
rect -4147 37 -4113 71
rect -4029 37 -3995 71
rect -3911 37 -3877 71
rect -3793 37 -3759 71
rect -3675 37 -3641 71
rect -3557 37 -3523 71
rect -3439 37 -3405 71
rect -3321 37 -3287 71
rect -3203 37 -3169 71
rect -3085 37 -3051 71
rect -2967 37 -2933 71
rect -2849 37 -2815 71
rect -2731 37 -2697 71
rect -2613 37 -2579 71
rect -2495 37 -2461 71
rect -2377 37 -2343 71
rect -2259 37 -2225 71
rect -2141 37 -2107 71
rect -2023 37 -1989 71
rect -1905 37 -1871 71
rect -1787 37 -1753 71
rect -1669 37 -1635 71
rect -1551 37 -1517 71
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect 1517 37 1551 71
rect 1635 37 1669 71
rect 1753 37 1787 71
rect 1871 37 1905 71
rect 1989 37 2023 71
rect 2107 37 2141 71
rect 2225 37 2259 71
rect 2343 37 2377 71
rect 2461 37 2495 71
rect 2579 37 2613 71
rect 2697 37 2731 71
rect 2815 37 2849 71
rect 2933 37 2967 71
rect 3051 37 3085 71
rect 3169 37 3203 71
rect 3287 37 3321 71
rect 3405 37 3439 71
rect 3523 37 3557 71
rect 3641 37 3675 71
rect 3759 37 3793 71
rect 3877 37 3911 71
rect 3995 37 4029 71
rect 4113 37 4147 71
rect 4231 37 4265 71
rect 4349 37 4383 71
rect -4383 -71 -4349 -37
rect -4265 -71 -4231 -37
rect -4147 -71 -4113 -37
rect -4029 -71 -3995 -37
rect -3911 -71 -3877 -37
rect -3793 -71 -3759 -37
rect -3675 -71 -3641 -37
rect -3557 -71 -3523 -37
rect -3439 -71 -3405 -37
rect -3321 -71 -3287 -37
rect -3203 -71 -3169 -37
rect -3085 -71 -3051 -37
rect -2967 -71 -2933 -37
rect -2849 -71 -2815 -37
rect -2731 -71 -2697 -37
rect -2613 -71 -2579 -37
rect -2495 -71 -2461 -37
rect -2377 -71 -2343 -37
rect -2259 -71 -2225 -37
rect -2141 -71 -2107 -37
rect -2023 -71 -1989 -37
rect -1905 -71 -1871 -37
rect -1787 -71 -1753 -37
rect -1669 -71 -1635 -37
rect -1551 -71 -1517 -37
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
rect 1517 -71 1551 -37
rect 1635 -71 1669 -37
rect 1753 -71 1787 -37
rect 1871 -71 1905 -37
rect 1989 -71 2023 -37
rect 2107 -71 2141 -37
rect 2225 -71 2259 -37
rect 2343 -71 2377 -37
rect 2461 -71 2495 -37
rect 2579 -71 2613 -37
rect 2697 -71 2731 -37
rect 2815 -71 2849 -37
rect 2933 -71 2967 -37
rect 3051 -71 3085 -37
rect 3169 -71 3203 -37
rect 3287 -71 3321 -37
rect 3405 -71 3439 -37
rect 3523 -71 3557 -37
rect 3641 -71 3675 -37
rect 3759 -71 3793 -37
rect 3877 -71 3911 -37
rect 3995 -71 4029 -37
rect 4113 -71 4147 -37
rect 4231 -71 4265 -37
rect 4349 -71 4383 -37
rect -4442 -706 -4408 -130
rect -4324 -706 -4290 -130
rect -4206 -706 -4172 -130
rect -4088 -706 -4054 -130
rect -3970 -706 -3936 -130
rect -3852 -706 -3818 -130
rect -3734 -706 -3700 -130
rect -3616 -706 -3582 -130
rect -3498 -706 -3464 -130
rect -3380 -706 -3346 -130
rect -3262 -706 -3228 -130
rect -3144 -706 -3110 -130
rect -3026 -706 -2992 -130
rect -2908 -706 -2874 -130
rect -2790 -706 -2756 -130
rect -2672 -706 -2638 -130
rect -2554 -706 -2520 -130
rect -2436 -706 -2402 -130
rect -2318 -706 -2284 -130
rect -2200 -706 -2166 -130
rect -2082 -706 -2048 -130
rect -1964 -706 -1930 -130
rect -1846 -706 -1812 -130
rect -1728 -706 -1694 -130
rect -1610 -706 -1576 -130
rect -1492 -706 -1458 -130
rect -1374 -706 -1340 -130
rect -1256 -706 -1222 -130
rect -1138 -706 -1104 -130
rect -1020 -706 -986 -130
rect -902 -706 -868 -130
rect -784 -706 -750 -130
rect -666 -706 -632 -130
rect -548 -706 -514 -130
rect -430 -706 -396 -130
rect -312 -706 -278 -130
rect -194 -706 -160 -130
rect -76 -706 -42 -130
rect 42 -706 76 -130
rect 160 -706 194 -130
rect 278 -706 312 -130
rect 396 -706 430 -130
rect 514 -706 548 -130
rect 632 -706 666 -130
rect 750 -706 784 -130
rect 868 -706 902 -130
rect 986 -706 1020 -130
rect 1104 -706 1138 -130
rect 1222 -706 1256 -130
rect 1340 -706 1374 -130
rect 1458 -706 1492 -130
rect 1576 -706 1610 -130
rect 1694 -706 1728 -130
rect 1812 -706 1846 -130
rect 1930 -706 1964 -130
rect 2048 -706 2082 -130
rect 2166 -706 2200 -130
rect 2284 -706 2318 -130
rect 2402 -706 2436 -130
rect 2520 -706 2554 -130
rect 2638 -706 2672 -130
rect 2756 -706 2790 -130
rect 2874 -706 2908 -130
rect 2992 -706 3026 -130
rect 3110 -706 3144 -130
rect 3228 -706 3262 -130
rect 3346 -706 3380 -130
rect 3464 -706 3498 -130
rect 3582 -706 3616 -130
rect 3700 -706 3734 -130
rect 3818 -706 3852 -130
rect 3936 -706 3970 -130
rect 4054 -706 4088 -130
rect 4172 -706 4206 -130
rect 4290 -706 4324 -130
rect 4408 -706 4442 -130
rect -4383 -799 -4349 -765
rect -4265 -799 -4231 -765
rect -4147 -799 -4113 -765
rect -4029 -799 -3995 -765
rect -3911 -799 -3877 -765
rect -3793 -799 -3759 -765
rect -3675 -799 -3641 -765
rect -3557 -799 -3523 -765
rect -3439 -799 -3405 -765
rect -3321 -799 -3287 -765
rect -3203 -799 -3169 -765
rect -3085 -799 -3051 -765
rect -2967 -799 -2933 -765
rect -2849 -799 -2815 -765
rect -2731 -799 -2697 -765
rect -2613 -799 -2579 -765
rect -2495 -799 -2461 -765
rect -2377 -799 -2343 -765
rect -2259 -799 -2225 -765
rect -2141 -799 -2107 -765
rect -2023 -799 -1989 -765
rect -1905 -799 -1871 -765
rect -1787 -799 -1753 -765
rect -1669 -799 -1635 -765
rect -1551 -799 -1517 -765
rect -1433 -799 -1399 -765
rect -1315 -799 -1281 -765
rect -1197 -799 -1163 -765
rect -1079 -799 -1045 -765
rect -961 -799 -927 -765
rect -843 -799 -809 -765
rect -725 -799 -691 -765
rect -607 -799 -573 -765
rect -489 -799 -455 -765
rect -371 -799 -337 -765
rect -253 -799 -219 -765
rect -135 -799 -101 -765
rect -17 -799 17 -765
rect 101 -799 135 -765
rect 219 -799 253 -765
rect 337 -799 371 -765
rect 455 -799 489 -765
rect 573 -799 607 -765
rect 691 -799 725 -765
rect 809 -799 843 -765
rect 927 -799 961 -765
rect 1045 -799 1079 -765
rect 1163 -799 1197 -765
rect 1281 -799 1315 -765
rect 1399 -799 1433 -765
rect 1517 -799 1551 -765
rect 1635 -799 1669 -765
rect 1753 -799 1787 -765
rect 1871 -799 1905 -765
rect 1989 -799 2023 -765
rect 2107 -799 2141 -765
rect 2225 -799 2259 -765
rect 2343 -799 2377 -765
rect 2461 -799 2495 -765
rect 2579 -799 2613 -765
rect 2697 -799 2731 -765
rect 2815 -799 2849 -765
rect 2933 -799 2967 -765
rect 3051 -799 3085 -765
rect 3169 -799 3203 -765
rect 3287 -799 3321 -765
rect 3405 -799 3439 -765
rect 3523 -799 3557 -765
rect 3641 -799 3675 -765
rect 3759 -799 3793 -765
rect 3877 -799 3911 -765
rect 3995 -799 4029 -765
rect 4113 -799 4147 -765
rect 4231 -799 4265 -765
rect 4349 -799 4383 -765
<< metal1 >>
rect -4395 799 -4337 805
rect -4395 765 -4383 799
rect -4349 765 -4337 799
rect -4395 759 -4337 765
rect -4277 799 -4219 805
rect -4277 765 -4265 799
rect -4231 765 -4219 799
rect -4277 759 -4219 765
rect -4159 799 -4101 805
rect -4159 765 -4147 799
rect -4113 765 -4101 799
rect -4159 759 -4101 765
rect -4041 799 -3983 805
rect -4041 765 -4029 799
rect -3995 765 -3983 799
rect -4041 759 -3983 765
rect -3923 799 -3865 805
rect -3923 765 -3911 799
rect -3877 765 -3865 799
rect -3923 759 -3865 765
rect -3805 799 -3747 805
rect -3805 765 -3793 799
rect -3759 765 -3747 799
rect -3805 759 -3747 765
rect -3687 799 -3629 805
rect -3687 765 -3675 799
rect -3641 765 -3629 799
rect -3687 759 -3629 765
rect -3569 799 -3511 805
rect -3569 765 -3557 799
rect -3523 765 -3511 799
rect -3569 759 -3511 765
rect -3451 799 -3393 805
rect -3451 765 -3439 799
rect -3405 765 -3393 799
rect -3451 759 -3393 765
rect -3333 799 -3275 805
rect -3333 765 -3321 799
rect -3287 765 -3275 799
rect -3333 759 -3275 765
rect -3215 799 -3157 805
rect -3215 765 -3203 799
rect -3169 765 -3157 799
rect -3215 759 -3157 765
rect -3097 799 -3039 805
rect -3097 765 -3085 799
rect -3051 765 -3039 799
rect -3097 759 -3039 765
rect -2979 799 -2921 805
rect -2979 765 -2967 799
rect -2933 765 -2921 799
rect -2979 759 -2921 765
rect -2861 799 -2803 805
rect -2861 765 -2849 799
rect -2815 765 -2803 799
rect -2861 759 -2803 765
rect -2743 799 -2685 805
rect -2743 765 -2731 799
rect -2697 765 -2685 799
rect -2743 759 -2685 765
rect -2625 799 -2567 805
rect -2625 765 -2613 799
rect -2579 765 -2567 799
rect -2625 759 -2567 765
rect -2507 799 -2449 805
rect -2507 765 -2495 799
rect -2461 765 -2449 799
rect -2507 759 -2449 765
rect -2389 799 -2331 805
rect -2389 765 -2377 799
rect -2343 765 -2331 799
rect -2389 759 -2331 765
rect -2271 799 -2213 805
rect -2271 765 -2259 799
rect -2225 765 -2213 799
rect -2271 759 -2213 765
rect -2153 799 -2095 805
rect -2153 765 -2141 799
rect -2107 765 -2095 799
rect -2153 759 -2095 765
rect -2035 799 -1977 805
rect -2035 765 -2023 799
rect -1989 765 -1977 799
rect -2035 759 -1977 765
rect -1917 799 -1859 805
rect -1917 765 -1905 799
rect -1871 765 -1859 799
rect -1917 759 -1859 765
rect -1799 799 -1741 805
rect -1799 765 -1787 799
rect -1753 765 -1741 799
rect -1799 759 -1741 765
rect -1681 799 -1623 805
rect -1681 765 -1669 799
rect -1635 765 -1623 799
rect -1681 759 -1623 765
rect -1563 799 -1505 805
rect -1563 765 -1551 799
rect -1517 765 -1505 799
rect -1563 759 -1505 765
rect -1445 799 -1387 805
rect -1445 765 -1433 799
rect -1399 765 -1387 799
rect -1445 759 -1387 765
rect -1327 799 -1269 805
rect -1327 765 -1315 799
rect -1281 765 -1269 799
rect -1327 759 -1269 765
rect -1209 799 -1151 805
rect -1209 765 -1197 799
rect -1163 765 -1151 799
rect -1209 759 -1151 765
rect -1091 799 -1033 805
rect -1091 765 -1079 799
rect -1045 765 -1033 799
rect -1091 759 -1033 765
rect -973 799 -915 805
rect -973 765 -961 799
rect -927 765 -915 799
rect -973 759 -915 765
rect -855 799 -797 805
rect -855 765 -843 799
rect -809 765 -797 799
rect -855 759 -797 765
rect -737 799 -679 805
rect -737 765 -725 799
rect -691 765 -679 799
rect -737 759 -679 765
rect -619 799 -561 805
rect -619 765 -607 799
rect -573 765 -561 799
rect -619 759 -561 765
rect -501 799 -443 805
rect -501 765 -489 799
rect -455 765 -443 799
rect -501 759 -443 765
rect -383 799 -325 805
rect -383 765 -371 799
rect -337 765 -325 799
rect -383 759 -325 765
rect -265 799 -207 805
rect -265 765 -253 799
rect -219 765 -207 799
rect -265 759 -207 765
rect -147 799 -89 805
rect -147 765 -135 799
rect -101 765 -89 799
rect -147 759 -89 765
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect 89 799 147 805
rect 89 765 101 799
rect 135 765 147 799
rect 89 759 147 765
rect 207 799 265 805
rect 207 765 219 799
rect 253 765 265 799
rect 207 759 265 765
rect 325 799 383 805
rect 325 765 337 799
rect 371 765 383 799
rect 325 759 383 765
rect 443 799 501 805
rect 443 765 455 799
rect 489 765 501 799
rect 443 759 501 765
rect 561 799 619 805
rect 561 765 573 799
rect 607 765 619 799
rect 561 759 619 765
rect 679 799 737 805
rect 679 765 691 799
rect 725 765 737 799
rect 679 759 737 765
rect 797 799 855 805
rect 797 765 809 799
rect 843 765 855 799
rect 797 759 855 765
rect 915 799 973 805
rect 915 765 927 799
rect 961 765 973 799
rect 915 759 973 765
rect 1033 799 1091 805
rect 1033 765 1045 799
rect 1079 765 1091 799
rect 1033 759 1091 765
rect 1151 799 1209 805
rect 1151 765 1163 799
rect 1197 765 1209 799
rect 1151 759 1209 765
rect 1269 799 1327 805
rect 1269 765 1281 799
rect 1315 765 1327 799
rect 1269 759 1327 765
rect 1387 799 1445 805
rect 1387 765 1399 799
rect 1433 765 1445 799
rect 1387 759 1445 765
rect 1505 799 1563 805
rect 1505 765 1517 799
rect 1551 765 1563 799
rect 1505 759 1563 765
rect 1623 799 1681 805
rect 1623 765 1635 799
rect 1669 765 1681 799
rect 1623 759 1681 765
rect 1741 799 1799 805
rect 1741 765 1753 799
rect 1787 765 1799 799
rect 1741 759 1799 765
rect 1859 799 1917 805
rect 1859 765 1871 799
rect 1905 765 1917 799
rect 1859 759 1917 765
rect 1977 799 2035 805
rect 1977 765 1989 799
rect 2023 765 2035 799
rect 1977 759 2035 765
rect 2095 799 2153 805
rect 2095 765 2107 799
rect 2141 765 2153 799
rect 2095 759 2153 765
rect 2213 799 2271 805
rect 2213 765 2225 799
rect 2259 765 2271 799
rect 2213 759 2271 765
rect 2331 799 2389 805
rect 2331 765 2343 799
rect 2377 765 2389 799
rect 2331 759 2389 765
rect 2449 799 2507 805
rect 2449 765 2461 799
rect 2495 765 2507 799
rect 2449 759 2507 765
rect 2567 799 2625 805
rect 2567 765 2579 799
rect 2613 765 2625 799
rect 2567 759 2625 765
rect 2685 799 2743 805
rect 2685 765 2697 799
rect 2731 765 2743 799
rect 2685 759 2743 765
rect 2803 799 2861 805
rect 2803 765 2815 799
rect 2849 765 2861 799
rect 2803 759 2861 765
rect 2921 799 2979 805
rect 2921 765 2933 799
rect 2967 765 2979 799
rect 2921 759 2979 765
rect 3039 799 3097 805
rect 3039 765 3051 799
rect 3085 765 3097 799
rect 3039 759 3097 765
rect 3157 799 3215 805
rect 3157 765 3169 799
rect 3203 765 3215 799
rect 3157 759 3215 765
rect 3275 799 3333 805
rect 3275 765 3287 799
rect 3321 765 3333 799
rect 3275 759 3333 765
rect 3393 799 3451 805
rect 3393 765 3405 799
rect 3439 765 3451 799
rect 3393 759 3451 765
rect 3511 799 3569 805
rect 3511 765 3523 799
rect 3557 765 3569 799
rect 3511 759 3569 765
rect 3629 799 3687 805
rect 3629 765 3641 799
rect 3675 765 3687 799
rect 3629 759 3687 765
rect 3747 799 3805 805
rect 3747 765 3759 799
rect 3793 765 3805 799
rect 3747 759 3805 765
rect 3865 799 3923 805
rect 3865 765 3877 799
rect 3911 765 3923 799
rect 3865 759 3923 765
rect 3983 799 4041 805
rect 3983 765 3995 799
rect 4029 765 4041 799
rect 3983 759 4041 765
rect 4101 799 4159 805
rect 4101 765 4113 799
rect 4147 765 4159 799
rect 4101 759 4159 765
rect 4219 799 4277 805
rect 4219 765 4231 799
rect 4265 765 4277 799
rect 4219 759 4277 765
rect 4337 799 4395 805
rect 4337 765 4349 799
rect 4383 765 4395 799
rect 4337 759 4395 765
rect -4448 706 -4402 718
rect -4448 130 -4442 706
rect -4408 130 -4402 706
rect -4448 118 -4402 130
rect -4330 706 -4284 718
rect -4330 130 -4324 706
rect -4290 130 -4284 706
rect -4330 118 -4284 130
rect -4212 706 -4166 718
rect -4212 130 -4206 706
rect -4172 130 -4166 706
rect -4212 118 -4166 130
rect -4094 706 -4048 718
rect -4094 130 -4088 706
rect -4054 130 -4048 706
rect -4094 118 -4048 130
rect -3976 706 -3930 718
rect -3976 130 -3970 706
rect -3936 130 -3930 706
rect -3976 118 -3930 130
rect -3858 706 -3812 718
rect -3858 130 -3852 706
rect -3818 130 -3812 706
rect -3858 118 -3812 130
rect -3740 706 -3694 718
rect -3740 130 -3734 706
rect -3700 130 -3694 706
rect -3740 118 -3694 130
rect -3622 706 -3576 718
rect -3622 130 -3616 706
rect -3582 130 -3576 706
rect -3622 118 -3576 130
rect -3504 706 -3458 718
rect -3504 130 -3498 706
rect -3464 130 -3458 706
rect -3504 118 -3458 130
rect -3386 706 -3340 718
rect -3386 130 -3380 706
rect -3346 130 -3340 706
rect -3386 118 -3340 130
rect -3268 706 -3222 718
rect -3268 130 -3262 706
rect -3228 130 -3222 706
rect -3268 118 -3222 130
rect -3150 706 -3104 718
rect -3150 130 -3144 706
rect -3110 130 -3104 706
rect -3150 118 -3104 130
rect -3032 706 -2986 718
rect -3032 130 -3026 706
rect -2992 130 -2986 706
rect -3032 118 -2986 130
rect -2914 706 -2868 718
rect -2914 130 -2908 706
rect -2874 130 -2868 706
rect -2914 118 -2868 130
rect -2796 706 -2750 718
rect -2796 130 -2790 706
rect -2756 130 -2750 706
rect -2796 118 -2750 130
rect -2678 706 -2632 718
rect -2678 130 -2672 706
rect -2638 130 -2632 706
rect -2678 118 -2632 130
rect -2560 706 -2514 718
rect -2560 130 -2554 706
rect -2520 130 -2514 706
rect -2560 118 -2514 130
rect -2442 706 -2396 718
rect -2442 130 -2436 706
rect -2402 130 -2396 706
rect -2442 118 -2396 130
rect -2324 706 -2278 718
rect -2324 130 -2318 706
rect -2284 130 -2278 706
rect -2324 118 -2278 130
rect -2206 706 -2160 718
rect -2206 130 -2200 706
rect -2166 130 -2160 706
rect -2206 118 -2160 130
rect -2088 706 -2042 718
rect -2088 130 -2082 706
rect -2048 130 -2042 706
rect -2088 118 -2042 130
rect -1970 706 -1924 718
rect -1970 130 -1964 706
rect -1930 130 -1924 706
rect -1970 118 -1924 130
rect -1852 706 -1806 718
rect -1852 130 -1846 706
rect -1812 130 -1806 706
rect -1852 118 -1806 130
rect -1734 706 -1688 718
rect -1734 130 -1728 706
rect -1694 130 -1688 706
rect -1734 118 -1688 130
rect -1616 706 -1570 718
rect -1616 130 -1610 706
rect -1576 130 -1570 706
rect -1616 118 -1570 130
rect -1498 706 -1452 718
rect -1498 130 -1492 706
rect -1458 130 -1452 706
rect -1498 118 -1452 130
rect -1380 706 -1334 718
rect -1380 130 -1374 706
rect -1340 130 -1334 706
rect -1380 118 -1334 130
rect -1262 706 -1216 718
rect -1262 130 -1256 706
rect -1222 130 -1216 706
rect -1262 118 -1216 130
rect -1144 706 -1098 718
rect -1144 130 -1138 706
rect -1104 130 -1098 706
rect -1144 118 -1098 130
rect -1026 706 -980 718
rect -1026 130 -1020 706
rect -986 130 -980 706
rect -1026 118 -980 130
rect -908 706 -862 718
rect -908 130 -902 706
rect -868 130 -862 706
rect -908 118 -862 130
rect -790 706 -744 718
rect -790 130 -784 706
rect -750 130 -744 706
rect -790 118 -744 130
rect -672 706 -626 718
rect -672 130 -666 706
rect -632 130 -626 706
rect -672 118 -626 130
rect -554 706 -508 718
rect -554 130 -548 706
rect -514 130 -508 706
rect -554 118 -508 130
rect -436 706 -390 718
rect -436 130 -430 706
rect -396 130 -390 706
rect -436 118 -390 130
rect -318 706 -272 718
rect -318 130 -312 706
rect -278 130 -272 706
rect -318 118 -272 130
rect -200 706 -154 718
rect -200 130 -194 706
rect -160 130 -154 706
rect -200 118 -154 130
rect -82 706 -36 718
rect -82 130 -76 706
rect -42 130 -36 706
rect -82 118 -36 130
rect 36 706 82 718
rect 36 130 42 706
rect 76 130 82 706
rect 36 118 82 130
rect 154 706 200 718
rect 154 130 160 706
rect 194 130 200 706
rect 154 118 200 130
rect 272 706 318 718
rect 272 130 278 706
rect 312 130 318 706
rect 272 118 318 130
rect 390 706 436 718
rect 390 130 396 706
rect 430 130 436 706
rect 390 118 436 130
rect 508 706 554 718
rect 508 130 514 706
rect 548 130 554 706
rect 508 118 554 130
rect 626 706 672 718
rect 626 130 632 706
rect 666 130 672 706
rect 626 118 672 130
rect 744 706 790 718
rect 744 130 750 706
rect 784 130 790 706
rect 744 118 790 130
rect 862 706 908 718
rect 862 130 868 706
rect 902 130 908 706
rect 862 118 908 130
rect 980 706 1026 718
rect 980 130 986 706
rect 1020 130 1026 706
rect 980 118 1026 130
rect 1098 706 1144 718
rect 1098 130 1104 706
rect 1138 130 1144 706
rect 1098 118 1144 130
rect 1216 706 1262 718
rect 1216 130 1222 706
rect 1256 130 1262 706
rect 1216 118 1262 130
rect 1334 706 1380 718
rect 1334 130 1340 706
rect 1374 130 1380 706
rect 1334 118 1380 130
rect 1452 706 1498 718
rect 1452 130 1458 706
rect 1492 130 1498 706
rect 1452 118 1498 130
rect 1570 706 1616 718
rect 1570 130 1576 706
rect 1610 130 1616 706
rect 1570 118 1616 130
rect 1688 706 1734 718
rect 1688 130 1694 706
rect 1728 130 1734 706
rect 1688 118 1734 130
rect 1806 706 1852 718
rect 1806 130 1812 706
rect 1846 130 1852 706
rect 1806 118 1852 130
rect 1924 706 1970 718
rect 1924 130 1930 706
rect 1964 130 1970 706
rect 1924 118 1970 130
rect 2042 706 2088 718
rect 2042 130 2048 706
rect 2082 130 2088 706
rect 2042 118 2088 130
rect 2160 706 2206 718
rect 2160 130 2166 706
rect 2200 130 2206 706
rect 2160 118 2206 130
rect 2278 706 2324 718
rect 2278 130 2284 706
rect 2318 130 2324 706
rect 2278 118 2324 130
rect 2396 706 2442 718
rect 2396 130 2402 706
rect 2436 130 2442 706
rect 2396 118 2442 130
rect 2514 706 2560 718
rect 2514 130 2520 706
rect 2554 130 2560 706
rect 2514 118 2560 130
rect 2632 706 2678 718
rect 2632 130 2638 706
rect 2672 130 2678 706
rect 2632 118 2678 130
rect 2750 706 2796 718
rect 2750 130 2756 706
rect 2790 130 2796 706
rect 2750 118 2796 130
rect 2868 706 2914 718
rect 2868 130 2874 706
rect 2908 130 2914 706
rect 2868 118 2914 130
rect 2986 706 3032 718
rect 2986 130 2992 706
rect 3026 130 3032 706
rect 2986 118 3032 130
rect 3104 706 3150 718
rect 3104 130 3110 706
rect 3144 130 3150 706
rect 3104 118 3150 130
rect 3222 706 3268 718
rect 3222 130 3228 706
rect 3262 130 3268 706
rect 3222 118 3268 130
rect 3340 706 3386 718
rect 3340 130 3346 706
rect 3380 130 3386 706
rect 3340 118 3386 130
rect 3458 706 3504 718
rect 3458 130 3464 706
rect 3498 130 3504 706
rect 3458 118 3504 130
rect 3576 706 3622 718
rect 3576 130 3582 706
rect 3616 130 3622 706
rect 3576 118 3622 130
rect 3694 706 3740 718
rect 3694 130 3700 706
rect 3734 130 3740 706
rect 3694 118 3740 130
rect 3812 706 3858 718
rect 3812 130 3818 706
rect 3852 130 3858 706
rect 3812 118 3858 130
rect 3930 706 3976 718
rect 3930 130 3936 706
rect 3970 130 3976 706
rect 3930 118 3976 130
rect 4048 706 4094 718
rect 4048 130 4054 706
rect 4088 130 4094 706
rect 4048 118 4094 130
rect 4166 706 4212 718
rect 4166 130 4172 706
rect 4206 130 4212 706
rect 4166 118 4212 130
rect 4284 706 4330 718
rect 4284 130 4290 706
rect 4324 130 4330 706
rect 4284 118 4330 130
rect 4402 706 4448 718
rect 4402 130 4408 706
rect 4442 130 4448 706
rect 4402 118 4448 130
rect -4395 71 -4337 77
rect -4395 37 -4383 71
rect -4349 37 -4337 71
rect -4395 31 -4337 37
rect -4277 71 -4219 77
rect -4277 37 -4265 71
rect -4231 37 -4219 71
rect -4277 31 -4219 37
rect -4159 71 -4101 77
rect -4159 37 -4147 71
rect -4113 37 -4101 71
rect -4159 31 -4101 37
rect -4041 71 -3983 77
rect -4041 37 -4029 71
rect -3995 37 -3983 71
rect -4041 31 -3983 37
rect -3923 71 -3865 77
rect -3923 37 -3911 71
rect -3877 37 -3865 71
rect -3923 31 -3865 37
rect -3805 71 -3747 77
rect -3805 37 -3793 71
rect -3759 37 -3747 71
rect -3805 31 -3747 37
rect -3687 71 -3629 77
rect -3687 37 -3675 71
rect -3641 37 -3629 71
rect -3687 31 -3629 37
rect -3569 71 -3511 77
rect -3569 37 -3557 71
rect -3523 37 -3511 71
rect -3569 31 -3511 37
rect -3451 71 -3393 77
rect -3451 37 -3439 71
rect -3405 37 -3393 71
rect -3451 31 -3393 37
rect -3333 71 -3275 77
rect -3333 37 -3321 71
rect -3287 37 -3275 71
rect -3333 31 -3275 37
rect -3215 71 -3157 77
rect -3215 37 -3203 71
rect -3169 37 -3157 71
rect -3215 31 -3157 37
rect -3097 71 -3039 77
rect -3097 37 -3085 71
rect -3051 37 -3039 71
rect -3097 31 -3039 37
rect -2979 71 -2921 77
rect -2979 37 -2967 71
rect -2933 37 -2921 71
rect -2979 31 -2921 37
rect -2861 71 -2803 77
rect -2861 37 -2849 71
rect -2815 37 -2803 71
rect -2861 31 -2803 37
rect -2743 71 -2685 77
rect -2743 37 -2731 71
rect -2697 37 -2685 71
rect -2743 31 -2685 37
rect -2625 71 -2567 77
rect -2625 37 -2613 71
rect -2579 37 -2567 71
rect -2625 31 -2567 37
rect -2507 71 -2449 77
rect -2507 37 -2495 71
rect -2461 37 -2449 71
rect -2507 31 -2449 37
rect -2389 71 -2331 77
rect -2389 37 -2377 71
rect -2343 37 -2331 71
rect -2389 31 -2331 37
rect -2271 71 -2213 77
rect -2271 37 -2259 71
rect -2225 37 -2213 71
rect -2271 31 -2213 37
rect -2153 71 -2095 77
rect -2153 37 -2141 71
rect -2107 37 -2095 71
rect -2153 31 -2095 37
rect -2035 71 -1977 77
rect -2035 37 -2023 71
rect -1989 37 -1977 71
rect -2035 31 -1977 37
rect -1917 71 -1859 77
rect -1917 37 -1905 71
rect -1871 37 -1859 71
rect -1917 31 -1859 37
rect -1799 71 -1741 77
rect -1799 37 -1787 71
rect -1753 37 -1741 71
rect -1799 31 -1741 37
rect -1681 71 -1623 77
rect -1681 37 -1669 71
rect -1635 37 -1623 71
rect -1681 31 -1623 37
rect -1563 71 -1505 77
rect -1563 37 -1551 71
rect -1517 37 -1505 71
rect -1563 31 -1505 37
rect -1445 71 -1387 77
rect -1445 37 -1433 71
rect -1399 37 -1387 71
rect -1445 31 -1387 37
rect -1327 71 -1269 77
rect -1327 37 -1315 71
rect -1281 37 -1269 71
rect -1327 31 -1269 37
rect -1209 71 -1151 77
rect -1209 37 -1197 71
rect -1163 37 -1151 71
rect -1209 31 -1151 37
rect -1091 71 -1033 77
rect -1091 37 -1079 71
rect -1045 37 -1033 71
rect -1091 31 -1033 37
rect -973 71 -915 77
rect -973 37 -961 71
rect -927 37 -915 71
rect -973 31 -915 37
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect 915 71 973 77
rect 915 37 927 71
rect 961 37 973 71
rect 915 31 973 37
rect 1033 71 1091 77
rect 1033 37 1045 71
rect 1079 37 1091 71
rect 1033 31 1091 37
rect 1151 71 1209 77
rect 1151 37 1163 71
rect 1197 37 1209 71
rect 1151 31 1209 37
rect 1269 71 1327 77
rect 1269 37 1281 71
rect 1315 37 1327 71
rect 1269 31 1327 37
rect 1387 71 1445 77
rect 1387 37 1399 71
rect 1433 37 1445 71
rect 1387 31 1445 37
rect 1505 71 1563 77
rect 1505 37 1517 71
rect 1551 37 1563 71
rect 1505 31 1563 37
rect 1623 71 1681 77
rect 1623 37 1635 71
rect 1669 37 1681 71
rect 1623 31 1681 37
rect 1741 71 1799 77
rect 1741 37 1753 71
rect 1787 37 1799 71
rect 1741 31 1799 37
rect 1859 71 1917 77
rect 1859 37 1871 71
rect 1905 37 1917 71
rect 1859 31 1917 37
rect 1977 71 2035 77
rect 1977 37 1989 71
rect 2023 37 2035 71
rect 1977 31 2035 37
rect 2095 71 2153 77
rect 2095 37 2107 71
rect 2141 37 2153 71
rect 2095 31 2153 37
rect 2213 71 2271 77
rect 2213 37 2225 71
rect 2259 37 2271 71
rect 2213 31 2271 37
rect 2331 71 2389 77
rect 2331 37 2343 71
rect 2377 37 2389 71
rect 2331 31 2389 37
rect 2449 71 2507 77
rect 2449 37 2461 71
rect 2495 37 2507 71
rect 2449 31 2507 37
rect 2567 71 2625 77
rect 2567 37 2579 71
rect 2613 37 2625 71
rect 2567 31 2625 37
rect 2685 71 2743 77
rect 2685 37 2697 71
rect 2731 37 2743 71
rect 2685 31 2743 37
rect 2803 71 2861 77
rect 2803 37 2815 71
rect 2849 37 2861 71
rect 2803 31 2861 37
rect 2921 71 2979 77
rect 2921 37 2933 71
rect 2967 37 2979 71
rect 2921 31 2979 37
rect 3039 71 3097 77
rect 3039 37 3051 71
rect 3085 37 3097 71
rect 3039 31 3097 37
rect 3157 71 3215 77
rect 3157 37 3169 71
rect 3203 37 3215 71
rect 3157 31 3215 37
rect 3275 71 3333 77
rect 3275 37 3287 71
rect 3321 37 3333 71
rect 3275 31 3333 37
rect 3393 71 3451 77
rect 3393 37 3405 71
rect 3439 37 3451 71
rect 3393 31 3451 37
rect 3511 71 3569 77
rect 3511 37 3523 71
rect 3557 37 3569 71
rect 3511 31 3569 37
rect 3629 71 3687 77
rect 3629 37 3641 71
rect 3675 37 3687 71
rect 3629 31 3687 37
rect 3747 71 3805 77
rect 3747 37 3759 71
rect 3793 37 3805 71
rect 3747 31 3805 37
rect 3865 71 3923 77
rect 3865 37 3877 71
rect 3911 37 3923 71
rect 3865 31 3923 37
rect 3983 71 4041 77
rect 3983 37 3995 71
rect 4029 37 4041 71
rect 3983 31 4041 37
rect 4101 71 4159 77
rect 4101 37 4113 71
rect 4147 37 4159 71
rect 4101 31 4159 37
rect 4219 71 4277 77
rect 4219 37 4231 71
rect 4265 37 4277 71
rect 4219 31 4277 37
rect 4337 71 4395 77
rect 4337 37 4349 71
rect 4383 37 4395 71
rect 4337 31 4395 37
rect -4395 -37 -4337 -31
rect -4395 -71 -4383 -37
rect -4349 -71 -4337 -37
rect -4395 -77 -4337 -71
rect -4277 -37 -4219 -31
rect -4277 -71 -4265 -37
rect -4231 -71 -4219 -37
rect -4277 -77 -4219 -71
rect -4159 -37 -4101 -31
rect -4159 -71 -4147 -37
rect -4113 -71 -4101 -37
rect -4159 -77 -4101 -71
rect -4041 -37 -3983 -31
rect -4041 -71 -4029 -37
rect -3995 -71 -3983 -37
rect -4041 -77 -3983 -71
rect -3923 -37 -3865 -31
rect -3923 -71 -3911 -37
rect -3877 -71 -3865 -37
rect -3923 -77 -3865 -71
rect -3805 -37 -3747 -31
rect -3805 -71 -3793 -37
rect -3759 -71 -3747 -37
rect -3805 -77 -3747 -71
rect -3687 -37 -3629 -31
rect -3687 -71 -3675 -37
rect -3641 -71 -3629 -37
rect -3687 -77 -3629 -71
rect -3569 -37 -3511 -31
rect -3569 -71 -3557 -37
rect -3523 -71 -3511 -37
rect -3569 -77 -3511 -71
rect -3451 -37 -3393 -31
rect -3451 -71 -3439 -37
rect -3405 -71 -3393 -37
rect -3451 -77 -3393 -71
rect -3333 -37 -3275 -31
rect -3333 -71 -3321 -37
rect -3287 -71 -3275 -37
rect -3333 -77 -3275 -71
rect -3215 -37 -3157 -31
rect -3215 -71 -3203 -37
rect -3169 -71 -3157 -37
rect -3215 -77 -3157 -71
rect -3097 -37 -3039 -31
rect -3097 -71 -3085 -37
rect -3051 -71 -3039 -37
rect -3097 -77 -3039 -71
rect -2979 -37 -2921 -31
rect -2979 -71 -2967 -37
rect -2933 -71 -2921 -37
rect -2979 -77 -2921 -71
rect -2861 -37 -2803 -31
rect -2861 -71 -2849 -37
rect -2815 -71 -2803 -37
rect -2861 -77 -2803 -71
rect -2743 -37 -2685 -31
rect -2743 -71 -2731 -37
rect -2697 -71 -2685 -37
rect -2743 -77 -2685 -71
rect -2625 -37 -2567 -31
rect -2625 -71 -2613 -37
rect -2579 -71 -2567 -37
rect -2625 -77 -2567 -71
rect -2507 -37 -2449 -31
rect -2507 -71 -2495 -37
rect -2461 -71 -2449 -37
rect -2507 -77 -2449 -71
rect -2389 -37 -2331 -31
rect -2389 -71 -2377 -37
rect -2343 -71 -2331 -37
rect -2389 -77 -2331 -71
rect -2271 -37 -2213 -31
rect -2271 -71 -2259 -37
rect -2225 -71 -2213 -37
rect -2271 -77 -2213 -71
rect -2153 -37 -2095 -31
rect -2153 -71 -2141 -37
rect -2107 -71 -2095 -37
rect -2153 -77 -2095 -71
rect -2035 -37 -1977 -31
rect -2035 -71 -2023 -37
rect -1989 -71 -1977 -37
rect -2035 -77 -1977 -71
rect -1917 -37 -1859 -31
rect -1917 -71 -1905 -37
rect -1871 -71 -1859 -37
rect -1917 -77 -1859 -71
rect -1799 -37 -1741 -31
rect -1799 -71 -1787 -37
rect -1753 -71 -1741 -37
rect -1799 -77 -1741 -71
rect -1681 -37 -1623 -31
rect -1681 -71 -1669 -37
rect -1635 -71 -1623 -37
rect -1681 -77 -1623 -71
rect -1563 -37 -1505 -31
rect -1563 -71 -1551 -37
rect -1517 -71 -1505 -37
rect -1563 -77 -1505 -71
rect -1445 -37 -1387 -31
rect -1445 -71 -1433 -37
rect -1399 -71 -1387 -37
rect -1445 -77 -1387 -71
rect -1327 -37 -1269 -31
rect -1327 -71 -1315 -37
rect -1281 -71 -1269 -37
rect -1327 -77 -1269 -71
rect -1209 -37 -1151 -31
rect -1209 -71 -1197 -37
rect -1163 -71 -1151 -37
rect -1209 -77 -1151 -71
rect -1091 -37 -1033 -31
rect -1091 -71 -1079 -37
rect -1045 -71 -1033 -37
rect -1091 -77 -1033 -71
rect -973 -37 -915 -31
rect -973 -71 -961 -37
rect -927 -71 -915 -37
rect -973 -77 -915 -71
rect -855 -37 -797 -31
rect -855 -71 -843 -37
rect -809 -71 -797 -37
rect -855 -77 -797 -71
rect -737 -37 -679 -31
rect -737 -71 -725 -37
rect -691 -71 -679 -37
rect -737 -77 -679 -71
rect -619 -37 -561 -31
rect -619 -71 -607 -37
rect -573 -71 -561 -37
rect -619 -77 -561 -71
rect -501 -37 -443 -31
rect -501 -71 -489 -37
rect -455 -71 -443 -37
rect -501 -77 -443 -71
rect -383 -37 -325 -31
rect -383 -71 -371 -37
rect -337 -71 -325 -37
rect -383 -77 -325 -71
rect -265 -37 -207 -31
rect -265 -71 -253 -37
rect -219 -71 -207 -37
rect -265 -77 -207 -71
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect 207 -37 265 -31
rect 207 -71 219 -37
rect 253 -71 265 -37
rect 207 -77 265 -71
rect 325 -37 383 -31
rect 325 -71 337 -37
rect 371 -71 383 -37
rect 325 -77 383 -71
rect 443 -37 501 -31
rect 443 -71 455 -37
rect 489 -71 501 -37
rect 443 -77 501 -71
rect 561 -37 619 -31
rect 561 -71 573 -37
rect 607 -71 619 -37
rect 561 -77 619 -71
rect 679 -37 737 -31
rect 679 -71 691 -37
rect 725 -71 737 -37
rect 679 -77 737 -71
rect 797 -37 855 -31
rect 797 -71 809 -37
rect 843 -71 855 -37
rect 797 -77 855 -71
rect 915 -37 973 -31
rect 915 -71 927 -37
rect 961 -71 973 -37
rect 915 -77 973 -71
rect 1033 -37 1091 -31
rect 1033 -71 1045 -37
rect 1079 -71 1091 -37
rect 1033 -77 1091 -71
rect 1151 -37 1209 -31
rect 1151 -71 1163 -37
rect 1197 -71 1209 -37
rect 1151 -77 1209 -71
rect 1269 -37 1327 -31
rect 1269 -71 1281 -37
rect 1315 -71 1327 -37
rect 1269 -77 1327 -71
rect 1387 -37 1445 -31
rect 1387 -71 1399 -37
rect 1433 -71 1445 -37
rect 1387 -77 1445 -71
rect 1505 -37 1563 -31
rect 1505 -71 1517 -37
rect 1551 -71 1563 -37
rect 1505 -77 1563 -71
rect 1623 -37 1681 -31
rect 1623 -71 1635 -37
rect 1669 -71 1681 -37
rect 1623 -77 1681 -71
rect 1741 -37 1799 -31
rect 1741 -71 1753 -37
rect 1787 -71 1799 -37
rect 1741 -77 1799 -71
rect 1859 -37 1917 -31
rect 1859 -71 1871 -37
rect 1905 -71 1917 -37
rect 1859 -77 1917 -71
rect 1977 -37 2035 -31
rect 1977 -71 1989 -37
rect 2023 -71 2035 -37
rect 1977 -77 2035 -71
rect 2095 -37 2153 -31
rect 2095 -71 2107 -37
rect 2141 -71 2153 -37
rect 2095 -77 2153 -71
rect 2213 -37 2271 -31
rect 2213 -71 2225 -37
rect 2259 -71 2271 -37
rect 2213 -77 2271 -71
rect 2331 -37 2389 -31
rect 2331 -71 2343 -37
rect 2377 -71 2389 -37
rect 2331 -77 2389 -71
rect 2449 -37 2507 -31
rect 2449 -71 2461 -37
rect 2495 -71 2507 -37
rect 2449 -77 2507 -71
rect 2567 -37 2625 -31
rect 2567 -71 2579 -37
rect 2613 -71 2625 -37
rect 2567 -77 2625 -71
rect 2685 -37 2743 -31
rect 2685 -71 2697 -37
rect 2731 -71 2743 -37
rect 2685 -77 2743 -71
rect 2803 -37 2861 -31
rect 2803 -71 2815 -37
rect 2849 -71 2861 -37
rect 2803 -77 2861 -71
rect 2921 -37 2979 -31
rect 2921 -71 2933 -37
rect 2967 -71 2979 -37
rect 2921 -77 2979 -71
rect 3039 -37 3097 -31
rect 3039 -71 3051 -37
rect 3085 -71 3097 -37
rect 3039 -77 3097 -71
rect 3157 -37 3215 -31
rect 3157 -71 3169 -37
rect 3203 -71 3215 -37
rect 3157 -77 3215 -71
rect 3275 -37 3333 -31
rect 3275 -71 3287 -37
rect 3321 -71 3333 -37
rect 3275 -77 3333 -71
rect 3393 -37 3451 -31
rect 3393 -71 3405 -37
rect 3439 -71 3451 -37
rect 3393 -77 3451 -71
rect 3511 -37 3569 -31
rect 3511 -71 3523 -37
rect 3557 -71 3569 -37
rect 3511 -77 3569 -71
rect 3629 -37 3687 -31
rect 3629 -71 3641 -37
rect 3675 -71 3687 -37
rect 3629 -77 3687 -71
rect 3747 -37 3805 -31
rect 3747 -71 3759 -37
rect 3793 -71 3805 -37
rect 3747 -77 3805 -71
rect 3865 -37 3923 -31
rect 3865 -71 3877 -37
rect 3911 -71 3923 -37
rect 3865 -77 3923 -71
rect 3983 -37 4041 -31
rect 3983 -71 3995 -37
rect 4029 -71 4041 -37
rect 3983 -77 4041 -71
rect 4101 -37 4159 -31
rect 4101 -71 4113 -37
rect 4147 -71 4159 -37
rect 4101 -77 4159 -71
rect 4219 -37 4277 -31
rect 4219 -71 4231 -37
rect 4265 -71 4277 -37
rect 4219 -77 4277 -71
rect 4337 -37 4395 -31
rect 4337 -71 4349 -37
rect 4383 -71 4395 -37
rect 4337 -77 4395 -71
rect -4448 -130 -4402 -118
rect -4448 -706 -4442 -130
rect -4408 -706 -4402 -130
rect -4448 -718 -4402 -706
rect -4330 -130 -4284 -118
rect -4330 -706 -4324 -130
rect -4290 -706 -4284 -130
rect -4330 -718 -4284 -706
rect -4212 -130 -4166 -118
rect -4212 -706 -4206 -130
rect -4172 -706 -4166 -130
rect -4212 -718 -4166 -706
rect -4094 -130 -4048 -118
rect -4094 -706 -4088 -130
rect -4054 -706 -4048 -130
rect -4094 -718 -4048 -706
rect -3976 -130 -3930 -118
rect -3976 -706 -3970 -130
rect -3936 -706 -3930 -130
rect -3976 -718 -3930 -706
rect -3858 -130 -3812 -118
rect -3858 -706 -3852 -130
rect -3818 -706 -3812 -130
rect -3858 -718 -3812 -706
rect -3740 -130 -3694 -118
rect -3740 -706 -3734 -130
rect -3700 -706 -3694 -130
rect -3740 -718 -3694 -706
rect -3622 -130 -3576 -118
rect -3622 -706 -3616 -130
rect -3582 -706 -3576 -130
rect -3622 -718 -3576 -706
rect -3504 -130 -3458 -118
rect -3504 -706 -3498 -130
rect -3464 -706 -3458 -130
rect -3504 -718 -3458 -706
rect -3386 -130 -3340 -118
rect -3386 -706 -3380 -130
rect -3346 -706 -3340 -130
rect -3386 -718 -3340 -706
rect -3268 -130 -3222 -118
rect -3268 -706 -3262 -130
rect -3228 -706 -3222 -130
rect -3268 -718 -3222 -706
rect -3150 -130 -3104 -118
rect -3150 -706 -3144 -130
rect -3110 -706 -3104 -130
rect -3150 -718 -3104 -706
rect -3032 -130 -2986 -118
rect -3032 -706 -3026 -130
rect -2992 -706 -2986 -130
rect -3032 -718 -2986 -706
rect -2914 -130 -2868 -118
rect -2914 -706 -2908 -130
rect -2874 -706 -2868 -130
rect -2914 -718 -2868 -706
rect -2796 -130 -2750 -118
rect -2796 -706 -2790 -130
rect -2756 -706 -2750 -130
rect -2796 -718 -2750 -706
rect -2678 -130 -2632 -118
rect -2678 -706 -2672 -130
rect -2638 -706 -2632 -130
rect -2678 -718 -2632 -706
rect -2560 -130 -2514 -118
rect -2560 -706 -2554 -130
rect -2520 -706 -2514 -130
rect -2560 -718 -2514 -706
rect -2442 -130 -2396 -118
rect -2442 -706 -2436 -130
rect -2402 -706 -2396 -130
rect -2442 -718 -2396 -706
rect -2324 -130 -2278 -118
rect -2324 -706 -2318 -130
rect -2284 -706 -2278 -130
rect -2324 -718 -2278 -706
rect -2206 -130 -2160 -118
rect -2206 -706 -2200 -130
rect -2166 -706 -2160 -130
rect -2206 -718 -2160 -706
rect -2088 -130 -2042 -118
rect -2088 -706 -2082 -130
rect -2048 -706 -2042 -130
rect -2088 -718 -2042 -706
rect -1970 -130 -1924 -118
rect -1970 -706 -1964 -130
rect -1930 -706 -1924 -130
rect -1970 -718 -1924 -706
rect -1852 -130 -1806 -118
rect -1852 -706 -1846 -130
rect -1812 -706 -1806 -130
rect -1852 -718 -1806 -706
rect -1734 -130 -1688 -118
rect -1734 -706 -1728 -130
rect -1694 -706 -1688 -130
rect -1734 -718 -1688 -706
rect -1616 -130 -1570 -118
rect -1616 -706 -1610 -130
rect -1576 -706 -1570 -130
rect -1616 -718 -1570 -706
rect -1498 -130 -1452 -118
rect -1498 -706 -1492 -130
rect -1458 -706 -1452 -130
rect -1498 -718 -1452 -706
rect -1380 -130 -1334 -118
rect -1380 -706 -1374 -130
rect -1340 -706 -1334 -130
rect -1380 -718 -1334 -706
rect -1262 -130 -1216 -118
rect -1262 -706 -1256 -130
rect -1222 -706 -1216 -130
rect -1262 -718 -1216 -706
rect -1144 -130 -1098 -118
rect -1144 -706 -1138 -130
rect -1104 -706 -1098 -130
rect -1144 -718 -1098 -706
rect -1026 -130 -980 -118
rect -1026 -706 -1020 -130
rect -986 -706 -980 -130
rect -1026 -718 -980 -706
rect -908 -130 -862 -118
rect -908 -706 -902 -130
rect -868 -706 -862 -130
rect -908 -718 -862 -706
rect -790 -130 -744 -118
rect -790 -706 -784 -130
rect -750 -706 -744 -130
rect -790 -718 -744 -706
rect -672 -130 -626 -118
rect -672 -706 -666 -130
rect -632 -706 -626 -130
rect -672 -718 -626 -706
rect -554 -130 -508 -118
rect -554 -706 -548 -130
rect -514 -706 -508 -130
rect -554 -718 -508 -706
rect -436 -130 -390 -118
rect -436 -706 -430 -130
rect -396 -706 -390 -130
rect -436 -718 -390 -706
rect -318 -130 -272 -118
rect -318 -706 -312 -130
rect -278 -706 -272 -130
rect -318 -718 -272 -706
rect -200 -130 -154 -118
rect -200 -706 -194 -130
rect -160 -706 -154 -130
rect -200 -718 -154 -706
rect -82 -130 -36 -118
rect -82 -706 -76 -130
rect -42 -706 -36 -130
rect -82 -718 -36 -706
rect 36 -130 82 -118
rect 36 -706 42 -130
rect 76 -706 82 -130
rect 36 -718 82 -706
rect 154 -130 200 -118
rect 154 -706 160 -130
rect 194 -706 200 -130
rect 154 -718 200 -706
rect 272 -130 318 -118
rect 272 -706 278 -130
rect 312 -706 318 -130
rect 272 -718 318 -706
rect 390 -130 436 -118
rect 390 -706 396 -130
rect 430 -706 436 -130
rect 390 -718 436 -706
rect 508 -130 554 -118
rect 508 -706 514 -130
rect 548 -706 554 -130
rect 508 -718 554 -706
rect 626 -130 672 -118
rect 626 -706 632 -130
rect 666 -706 672 -130
rect 626 -718 672 -706
rect 744 -130 790 -118
rect 744 -706 750 -130
rect 784 -706 790 -130
rect 744 -718 790 -706
rect 862 -130 908 -118
rect 862 -706 868 -130
rect 902 -706 908 -130
rect 862 -718 908 -706
rect 980 -130 1026 -118
rect 980 -706 986 -130
rect 1020 -706 1026 -130
rect 980 -718 1026 -706
rect 1098 -130 1144 -118
rect 1098 -706 1104 -130
rect 1138 -706 1144 -130
rect 1098 -718 1144 -706
rect 1216 -130 1262 -118
rect 1216 -706 1222 -130
rect 1256 -706 1262 -130
rect 1216 -718 1262 -706
rect 1334 -130 1380 -118
rect 1334 -706 1340 -130
rect 1374 -706 1380 -130
rect 1334 -718 1380 -706
rect 1452 -130 1498 -118
rect 1452 -706 1458 -130
rect 1492 -706 1498 -130
rect 1452 -718 1498 -706
rect 1570 -130 1616 -118
rect 1570 -706 1576 -130
rect 1610 -706 1616 -130
rect 1570 -718 1616 -706
rect 1688 -130 1734 -118
rect 1688 -706 1694 -130
rect 1728 -706 1734 -130
rect 1688 -718 1734 -706
rect 1806 -130 1852 -118
rect 1806 -706 1812 -130
rect 1846 -706 1852 -130
rect 1806 -718 1852 -706
rect 1924 -130 1970 -118
rect 1924 -706 1930 -130
rect 1964 -706 1970 -130
rect 1924 -718 1970 -706
rect 2042 -130 2088 -118
rect 2042 -706 2048 -130
rect 2082 -706 2088 -130
rect 2042 -718 2088 -706
rect 2160 -130 2206 -118
rect 2160 -706 2166 -130
rect 2200 -706 2206 -130
rect 2160 -718 2206 -706
rect 2278 -130 2324 -118
rect 2278 -706 2284 -130
rect 2318 -706 2324 -130
rect 2278 -718 2324 -706
rect 2396 -130 2442 -118
rect 2396 -706 2402 -130
rect 2436 -706 2442 -130
rect 2396 -718 2442 -706
rect 2514 -130 2560 -118
rect 2514 -706 2520 -130
rect 2554 -706 2560 -130
rect 2514 -718 2560 -706
rect 2632 -130 2678 -118
rect 2632 -706 2638 -130
rect 2672 -706 2678 -130
rect 2632 -718 2678 -706
rect 2750 -130 2796 -118
rect 2750 -706 2756 -130
rect 2790 -706 2796 -130
rect 2750 -718 2796 -706
rect 2868 -130 2914 -118
rect 2868 -706 2874 -130
rect 2908 -706 2914 -130
rect 2868 -718 2914 -706
rect 2986 -130 3032 -118
rect 2986 -706 2992 -130
rect 3026 -706 3032 -130
rect 2986 -718 3032 -706
rect 3104 -130 3150 -118
rect 3104 -706 3110 -130
rect 3144 -706 3150 -130
rect 3104 -718 3150 -706
rect 3222 -130 3268 -118
rect 3222 -706 3228 -130
rect 3262 -706 3268 -130
rect 3222 -718 3268 -706
rect 3340 -130 3386 -118
rect 3340 -706 3346 -130
rect 3380 -706 3386 -130
rect 3340 -718 3386 -706
rect 3458 -130 3504 -118
rect 3458 -706 3464 -130
rect 3498 -706 3504 -130
rect 3458 -718 3504 -706
rect 3576 -130 3622 -118
rect 3576 -706 3582 -130
rect 3616 -706 3622 -130
rect 3576 -718 3622 -706
rect 3694 -130 3740 -118
rect 3694 -706 3700 -130
rect 3734 -706 3740 -130
rect 3694 -718 3740 -706
rect 3812 -130 3858 -118
rect 3812 -706 3818 -130
rect 3852 -706 3858 -130
rect 3812 -718 3858 -706
rect 3930 -130 3976 -118
rect 3930 -706 3936 -130
rect 3970 -706 3976 -130
rect 3930 -718 3976 -706
rect 4048 -130 4094 -118
rect 4048 -706 4054 -130
rect 4088 -706 4094 -130
rect 4048 -718 4094 -706
rect 4166 -130 4212 -118
rect 4166 -706 4172 -130
rect 4206 -706 4212 -130
rect 4166 -718 4212 -706
rect 4284 -130 4330 -118
rect 4284 -706 4290 -130
rect 4324 -706 4330 -130
rect 4284 -718 4330 -706
rect 4402 -130 4448 -118
rect 4402 -706 4408 -130
rect 4442 -706 4448 -130
rect 4402 -718 4448 -706
rect -4395 -765 -4337 -759
rect -4395 -799 -4383 -765
rect -4349 -799 -4337 -765
rect -4395 -805 -4337 -799
rect -4277 -765 -4219 -759
rect -4277 -799 -4265 -765
rect -4231 -799 -4219 -765
rect -4277 -805 -4219 -799
rect -4159 -765 -4101 -759
rect -4159 -799 -4147 -765
rect -4113 -799 -4101 -765
rect -4159 -805 -4101 -799
rect -4041 -765 -3983 -759
rect -4041 -799 -4029 -765
rect -3995 -799 -3983 -765
rect -4041 -805 -3983 -799
rect -3923 -765 -3865 -759
rect -3923 -799 -3911 -765
rect -3877 -799 -3865 -765
rect -3923 -805 -3865 -799
rect -3805 -765 -3747 -759
rect -3805 -799 -3793 -765
rect -3759 -799 -3747 -765
rect -3805 -805 -3747 -799
rect -3687 -765 -3629 -759
rect -3687 -799 -3675 -765
rect -3641 -799 -3629 -765
rect -3687 -805 -3629 -799
rect -3569 -765 -3511 -759
rect -3569 -799 -3557 -765
rect -3523 -799 -3511 -765
rect -3569 -805 -3511 -799
rect -3451 -765 -3393 -759
rect -3451 -799 -3439 -765
rect -3405 -799 -3393 -765
rect -3451 -805 -3393 -799
rect -3333 -765 -3275 -759
rect -3333 -799 -3321 -765
rect -3287 -799 -3275 -765
rect -3333 -805 -3275 -799
rect -3215 -765 -3157 -759
rect -3215 -799 -3203 -765
rect -3169 -799 -3157 -765
rect -3215 -805 -3157 -799
rect -3097 -765 -3039 -759
rect -3097 -799 -3085 -765
rect -3051 -799 -3039 -765
rect -3097 -805 -3039 -799
rect -2979 -765 -2921 -759
rect -2979 -799 -2967 -765
rect -2933 -799 -2921 -765
rect -2979 -805 -2921 -799
rect -2861 -765 -2803 -759
rect -2861 -799 -2849 -765
rect -2815 -799 -2803 -765
rect -2861 -805 -2803 -799
rect -2743 -765 -2685 -759
rect -2743 -799 -2731 -765
rect -2697 -799 -2685 -765
rect -2743 -805 -2685 -799
rect -2625 -765 -2567 -759
rect -2625 -799 -2613 -765
rect -2579 -799 -2567 -765
rect -2625 -805 -2567 -799
rect -2507 -765 -2449 -759
rect -2507 -799 -2495 -765
rect -2461 -799 -2449 -765
rect -2507 -805 -2449 -799
rect -2389 -765 -2331 -759
rect -2389 -799 -2377 -765
rect -2343 -799 -2331 -765
rect -2389 -805 -2331 -799
rect -2271 -765 -2213 -759
rect -2271 -799 -2259 -765
rect -2225 -799 -2213 -765
rect -2271 -805 -2213 -799
rect -2153 -765 -2095 -759
rect -2153 -799 -2141 -765
rect -2107 -799 -2095 -765
rect -2153 -805 -2095 -799
rect -2035 -765 -1977 -759
rect -2035 -799 -2023 -765
rect -1989 -799 -1977 -765
rect -2035 -805 -1977 -799
rect -1917 -765 -1859 -759
rect -1917 -799 -1905 -765
rect -1871 -799 -1859 -765
rect -1917 -805 -1859 -799
rect -1799 -765 -1741 -759
rect -1799 -799 -1787 -765
rect -1753 -799 -1741 -765
rect -1799 -805 -1741 -799
rect -1681 -765 -1623 -759
rect -1681 -799 -1669 -765
rect -1635 -799 -1623 -765
rect -1681 -805 -1623 -799
rect -1563 -765 -1505 -759
rect -1563 -799 -1551 -765
rect -1517 -799 -1505 -765
rect -1563 -805 -1505 -799
rect -1445 -765 -1387 -759
rect -1445 -799 -1433 -765
rect -1399 -799 -1387 -765
rect -1445 -805 -1387 -799
rect -1327 -765 -1269 -759
rect -1327 -799 -1315 -765
rect -1281 -799 -1269 -765
rect -1327 -805 -1269 -799
rect -1209 -765 -1151 -759
rect -1209 -799 -1197 -765
rect -1163 -799 -1151 -765
rect -1209 -805 -1151 -799
rect -1091 -765 -1033 -759
rect -1091 -799 -1079 -765
rect -1045 -799 -1033 -765
rect -1091 -805 -1033 -799
rect -973 -765 -915 -759
rect -973 -799 -961 -765
rect -927 -799 -915 -765
rect -973 -805 -915 -799
rect -855 -765 -797 -759
rect -855 -799 -843 -765
rect -809 -799 -797 -765
rect -855 -805 -797 -799
rect -737 -765 -679 -759
rect -737 -799 -725 -765
rect -691 -799 -679 -765
rect -737 -805 -679 -799
rect -619 -765 -561 -759
rect -619 -799 -607 -765
rect -573 -799 -561 -765
rect -619 -805 -561 -799
rect -501 -765 -443 -759
rect -501 -799 -489 -765
rect -455 -799 -443 -765
rect -501 -805 -443 -799
rect -383 -765 -325 -759
rect -383 -799 -371 -765
rect -337 -799 -325 -765
rect -383 -805 -325 -799
rect -265 -765 -207 -759
rect -265 -799 -253 -765
rect -219 -799 -207 -765
rect -265 -805 -207 -799
rect -147 -765 -89 -759
rect -147 -799 -135 -765
rect -101 -799 -89 -765
rect -147 -805 -89 -799
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect 89 -765 147 -759
rect 89 -799 101 -765
rect 135 -799 147 -765
rect 89 -805 147 -799
rect 207 -765 265 -759
rect 207 -799 219 -765
rect 253 -799 265 -765
rect 207 -805 265 -799
rect 325 -765 383 -759
rect 325 -799 337 -765
rect 371 -799 383 -765
rect 325 -805 383 -799
rect 443 -765 501 -759
rect 443 -799 455 -765
rect 489 -799 501 -765
rect 443 -805 501 -799
rect 561 -765 619 -759
rect 561 -799 573 -765
rect 607 -799 619 -765
rect 561 -805 619 -799
rect 679 -765 737 -759
rect 679 -799 691 -765
rect 725 -799 737 -765
rect 679 -805 737 -799
rect 797 -765 855 -759
rect 797 -799 809 -765
rect 843 -799 855 -765
rect 797 -805 855 -799
rect 915 -765 973 -759
rect 915 -799 927 -765
rect 961 -799 973 -765
rect 915 -805 973 -799
rect 1033 -765 1091 -759
rect 1033 -799 1045 -765
rect 1079 -799 1091 -765
rect 1033 -805 1091 -799
rect 1151 -765 1209 -759
rect 1151 -799 1163 -765
rect 1197 -799 1209 -765
rect 1151 -805 1209 -799
rect 1269 -765 1327 -759
rect 1269 -799 1281 -765
rect 1315 -799 1327 -765
rect 1269 -805 1327 -799
rect 1387 -765 1445 -759
rect 1387 -799 1399 -765
rect 1433 -799 1445 -765
rect 1387 -805 1445 -799
rect 1505 -765 1563 -759
rect 1505 -799 1517 -765
rect 1551 -799 1563 -765
rect 1505 -805 1563 -799
rect 1623 -765 1681 -759
rect 1623 -799 1635 -765
rect 1669 -799 1681 -765
rect 1623 -805 1681 -799
rect 1741 -765 1799 -759
rect 1741 -799 1753 -765
rect 1787 -799 1799 -765
rect 1741 -805 1799 -799
rect 1859 -765 1917 -759
rect 1859 -799 1871 -765
rect 1905 -799 1917 -765
rect 1859 -805 1917 -799
rect 1977 -765 2035 -759
rect 1977 -799 1989 -765
rect 2023 -799 2035 -765
rect 1977 -805 2035 -799
rect 2095 -765 2153 -759
rect 2095 -799 2107 -765
rect 2141 -799 2153 -765
rect 2095 -805 2153 -799
rect 2213 -765 2271 -759
rect 2213 -799 2225 -765
rect 2259 -799 2271 -765
rect 2213 -805 2271 -799
rect 2331 -765 2389 -759
rect 2331 -799 2343 -765
rect 2377 -799 2389 -765
rect 2331 -805 2389 -799
rect 2449 -765 2507 -759
rect 2449 -799 2461 -765
rect 2495 -799 2507 -765
rect 2449 -805 2507 -799
rect 2567 -765 2625 -759
rect 2567 -799 2579 -765
rect 2613 -799 2625 -765
rect 2567 -805 2625 -799
rect 2685 -765 2743 -759
rect 2685 -799 2697 -765
rect 2731 -799 2743 -765
rect 2685 -805 2743 -799
rect 2803 -765 2861 -759
rect 2803 -799 2815 -765
rect 2849 -799 2861 -765
rect 2803 -805 2861 -799
rect 2921 -765 2979 -759
rect 2921 -799 2933 -765
rect 2967 -799 2979 -765
rect 2921 -805 2979 -799
rect 3039 -765 3097 -759
rect 3039 -799 3051 -765
rect 3085 -799 3097 -765
rect 3039 -805 3097 -799
rect 3157 -765 3215 -759
rect 3157 -799 3169 -765
rect 3203 -799 3215 -765
rect 3157 -805 3215 -799
rect 3275 -765 3333 -759
rect 3275 -799 3287 -765
rect 3321 -799 3333 -765
rect 3275 -805 3333 -799
rect 3393 -765 3451 -759
rect 3393 -799 3405 -765
rect 3439 -799 3451 -765
rect 3393 -805 3451 -799
rect 3511 -765 3569 -759
rect 3511 -799 3523 -765
rect 3557 -799 3569 -765
rect 3511 -805 3569 -799
rect 3629 -765 3687 -759
rect 3629 -799 3641 -765
rect 3675 -799 3687 -765
rect 3629 -805 3687 -799
rect 3747 -765 3805 -759
rect 3747 -799 3759 -765
rect 3793 -799 3805 -765
rect 3747 -805 3805 -799
rect 3865 -765 3923 -759
rect 3865 -799 3877 -765
rect 3911 -799 3923 -765
rect 3865 -805 3923 -799
rect 3983 -765 4041 -759
rect 3983 -799 3995 -765
rect 4029 -799 4041 -765
rect 3983 -805 4041 -799
rect 4101 -765 4159 -759
rect 4101 -799 4113 -765
rect 4147 -799 4159 -765
rect 4101 -805 4159 -799
rect 4219 -765 4277 -759
rect 4219 -799 4231 -765
rect 4265 -799 4277 -765
rect 4219 -805 4277 -799
rect 4337 -765 4395 -759
rect 4337 -799 4349 -765
rect 4383 -799 4395 -765
rect 4337 -805 4395 -799
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -4539 -884 4539 884
string parameters w 3 l 0.3 m 2 nf 75 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
